magic
tech sky130A
magscale 1 2
timestamp 1672336121
<< obsli1 >>
rect 1104 2159 569664 684369
<< obsm1 >>
rect 382 2128 570754 684400
<< metal2 >>
rect 8390 685869 8446 686669
rect 24214 685869 24270 686669
rect 40038 685869 40094 686669
rect 55862 685869 55918 686669
rect 71686 685869 71742 686669
rect 87510 685869 87566 686669
rect 103334 685869 103390 686669
rect 119158 685869 119214 686669
rect 134982 685869 135038 686669
rect 150806 685869 150862 686669
rect 166630 685869 166686 686669
rect 182454 685869 182510 686669
rect 198278 685869 198334 686669
rect 214102 685869 214158 686669
rect 229926 685869 229982 686669
rect 245750 685869 245806 686669
rect 261574 685869 261630 686669
rect 277398 685869 277454 686669
rect 293222 685869 293278 686669
rect 309046 685869 309102 686669
rect 324870 685869 324926 686669
rect 340694 685869 340750 686669
rect 356518 685869 356574 686669
rect 372342 685869 372398 686669
rect 388166 685869 388222 686669
rect 403990 685869 404046 686669
rect 419814 685869 419870 686669
rect 435638 685869 435694 686669
rect 451462 685869 451518 686669
rect 467286 685869 467342 686669
rect 483110 685869 483166 686669
rect 498934 685869 498990 686669
rect 514758 685869 514814 686669
rect 530582 685869 530638 686669
rect 546406 685869 546462 686669
rect 562230 685869 562286 686669
rect 13174 0 13230 800
rect 14278 0 14334 800
rect 15382 0 15438 800
rect 16486 0 16542 800
rect 17590 0 17646 800
rect 18694 0 18750 800
rect 19798 0 19854 800
rect 20902 0 20958 800
rect 22006 0 22062 800
rect 23110 0 23166 800
rect 24214 0 24270 800
rect 25318 0 25374 800
rect 26422 0 26478 800
rect 27526 0 27582 800
rect 28630 0 28686 800
rect 29734 0 29790 800
rect 30838 0 30894 800
rect 31942 0 31998 800
rect 33046 0 33102 800
rect 34150 0 34206 800
rect 35254 0 35310 800
rect 36358 0 36414 800
rect 37462 0 37518 800
rect 38566 0 38622 800
rect 39670 0 39726 800
rect 40774 0 40830 800
rect 41878 0 41934 800
rect 42982 0 43038 800
rect 44086 0 44142 800
rect 45190 0 45246 800
rect 46294 0 46350 800
rect 47398 0 47454 800
rect 48502 0 48558 800
rect 49606 0 49662 800
rect 50710 0 50766 800
rect 51814 0 51870 800
rect 52918 0 52974 800
rect 54022 0 54078 800
rect 55126 0 55182 800
rect 56230 0 56286 800
rect 57334 0 57390 800
rect 58438 0 58494 800
rect 59542 0 59598 800
rect 60646 0 60702 800
rect 61750 0 61806 800
rect 62854 0 62910 800
rect 63958 0 64014 800
rect 65062 0 65118 800
rect 66166 0 66222 800
rect 67270 0 67326 800
rect 68374 0 68430 800
rect 69478 0 69534 800
rect 70582 0 70638 800
rect 71686 0 71742 800
rect 72790 0 72846 800
rect 73894 0 73950 800
rect 74998 0 75054 800
rect 76102 0 76158 800
rect 77206 0 77262 800
rect 78310 0 78366 800
rect 79414 0 79470 800
rect 80518 0 80574 800
rect 81622 0 81678 800
rect 82726 0 82782 800
rect 83830 0 83886 800
rect 84934 0 84990 800
rect 86038 0 86094 800
rect 87142 0 87198 800
rect 88246 0 88302 800
rect 89350 0 89406 800
rect 90454 0 90510 800
rect 91558 0 91614 800
rect 92662 0 92718 800
rect 93766 0 93822 800
rect 94870 0 94926 800
rect 95974 0 96030 800
rect 97078 0 97134 800
rect 98182 0 98238 800
rect 99286 0 99342 800
rect 100390 0 100446 800
rect 101494 0 101550 800
rect 102598 0 102654 800
rect 103702 0 103758 800
rect 104806 0 104862 800
rect 105910 0 105966 800
rect 107014 0 107070 800
rect 108118 0 108174 800
rect 109222 0 109278 800
rect 110326 0 110382 800
rect 111430 0 111486 800
rect 112534 0 112590 800
rect 113638 0 113694 800
rect 114742 0 114798 800
rect 115846 0 115902 800
rect 116950 0 117006 800
rect 118054 0 118110 800
rect 119158 0 119214 800
rect 120262 0 120318 800
rect 121366 0 121422 800
rect 122470 0 122526 800
rect 123574 0 123630 800
rect 124678 0 124734 800
rect 125782 0 125838 800
rect 126886 0 126942 800
rect 127990 0 128046 800
rect 129094 0 129150 800
rect 130198 0 130254 800
rect 131302 0 131358 800
rect 132406 0 132462 800
rect 133510 0 133566 800
rect 134614 0 134670 800
rect 135718 0 135774 800
rect 136822 0 136878 800
rect 137926 0 137982 800
rect 139030 0 139086 800
rect 140134 0 140190 800
rect 141238 0 141294 800
rect 142342 0 142398 800
rect 143446 0 143502 800
rect 144550 0 144606 800
rect 145654 0 145710 800
rect 146758 0 146814 800
rect 147862 0 147918 800
rect 148966 0 149022 800
rect 150070 0 150126 800
rect 151174 0 151230 800
rect 152278 0 152334 800
rect 153382 0 153438 800
rect 154486 0 154542 800
rect 155590 0 155646 800
rect 156694 0 156750 800
rect 157798 0 157854 800
rect 158902 0 158958 800
rect 160006 0 160062 800
rect 161110 0 161166 800
rect 162214 0 162270 800
rect 163318 0 163374 800
rect 164422 0 164478 800
rect 165526 0 165582 800
rect 166630 0 166686 800
rect 167734 0 167790 800
rect 168838 0 168894 800
rect 169942 0 169998 800
rect 171046 0 171102 800
rect 172150 0 172206 800
rect 173254 0 173310 800
rect 174358 0 174414 800
rect 175462 0 175518 800
rect 176566 0 176622 800
rect 177670 0 177726 800
rect 178774 0 178830 800
rect 179878 0 179934 800
rect 180982 0 181038 800
rect 182086 0 182142 800
rect 183190 0 183246 800
rect 184294 0 184350 800
rect 185398 0 185454 800
rect 186502 0 186558 800
rect 187606 0 187662 800
rect 188710 0 188766 800
rect 189814 0 189870 800
rect 190918 0 190974 800
rect 192022 0 192078 800
rect 193126 0 193182 800
rect 194230 0 194286 800
rect 195334 0 195390 800
rect 196438 0 196494 800
rect 197542 0 197598 800
rect 198646 0 198702 800
rect 199750 0 199806 800
rect 200854 0 200910 800
rect 201958 0 202014 800
rect 203062 0 203118 800
rect 204166 0 204222 800
rect 205270 0 205326 800
rect 206374 0 206430 800
rect 207478 0 207534 800
rect 208582 0 208638 800
rect 209686 0 209742 800
rect 210790 0 210846 800
rect 211894 0 211950 800
rect 212998 0 213054 800
rect 214102 0 214158 800
rect 215206 0 215262 800
rect 216310 0 216366 800
rect 217414 0 217470 800
rect 218518 0 218574 800
rect 219622 0 219678 800
rect 220726 0 220782 800
rect 221830 0 221886 800
rect 222934 0 222990 800
rect 224038 0 224094 800
rect 225142 0 225198 800
rect 226246 0 226302 800
rect 227350 0 227406 800
rect 228454 0 228510 800
rect 229558 0 229614 800
rect 230662 0 230718 800
rect 231766 0 231822 800
rect 232870 0 232926 800
rect 233974 0 234030 800
rect 235078 0 235134 800
rect 236182 0 236238 800
rect 237286 0 237342 800
rect 238390 0 238446 800
rect 239494 0 239550 800
rect 240598 0 240654 800
rect 241702 0 241758 800
rect 242806 0 242862 800
rect 243910 0 243966 800
rect 245014 0 245070 800
rect 246118 0 246174 800
rect 247222 0 247278 800
rect 248326 0 248382 800
rect 249430 0 249486 800
rect 250534 0 250590 800
rect 251638 0 251694 800
rect 252742 0 252798 800
rect 253846 0 253902 800
rect 254950 0 255006 800
rect 256054 0 256110 800
rect 257158 0 257214 800
rect 258262 0 258318 800
rect 259366 0 259422 800
rect 260470 0 260526 800
rect 261574 0 261630 800
rect 262678 0 262734 800
rect 263782 0 263838 800
rect 264886 0 264942 800
rect 265990 0 266046 800
rect 267094 0 267150 800
rect 268198 0 268254 800
rect 269302 0 269358 800
rect 270406 0 270462 800
rect 271510 0 271566 800
rect 272614 0 272670 800
rect 273718 0 273774 800
rect 274822 0 274878 800
rect 275926 0 275982 800
rect 277030 0 277086 800
rect 278134 0 278190 800
rect 279238 0 279294 800
rect 280342 0 280398 800
rect 281446 0 281502 800
rect 282550 0 282606 800
rect 283654 0 283710 800
rect 284758 0 284814 800
rect 285862 0 285918 800
rect 286966 0 287022 800
rect 288070 0 288126 800
rect 289174 0 289230 800
rect 290278 0 290334 800
rect 291382 0 291438 800
rect 292486 0 292542 800
rect 293590 0 293646 800
rect 294694 0 294750 800
rect 295798 0 295854 800
rect 296902 0 296958 800
rect 298006 0 298062 800
rect 299110 0 299166 800
rect 300214 0 300270 800
rect 301318 0 301374 800
rect 302422 0 302478 800
rect 303526 0 303582 800
rect 304630 0 304686 800
rect 305734 0 305790 800
rect 306838 0 306894 800
rect 307942 0 307998 800
rect 309046 0 309102 800
rect 310150 0 310206 800
rect 311254 0 311310 800
rect 312358 0 312414 800
rect 313462 0 313518 800
rect 314566 0 314622 800
rect 315670 0 315726 800
rect 316774 0 316830 800
rect 317878 0 317934 800
rect 318982 0 319038 800
rect 320086 0 320142 800
rect 321190 0 321246 800
rect 322294 0 322350 800
rect 323398 0 323454 800
rect 324502 0 324558 800
rect 325606 0 325662 800
rect 326710 0 326766 800
rect 327814 0 327870 800
rect 328918 0 328974 800
rect 330022 0 330078 800
rect 331126 0 331182 800
rect 332230 0 332286 800
rect 333334 0 333390 800
rect 334438 0 334494 800
rect 335542 0 335598 800
rect 336646 0 336702 800
rect 337750 0 337806 800
rect 338854 0 338910 800
rect 339958 0 340014 800
rect 341062 0 341118 800
rect 342166 0 342222 800
rect 343270 0 343326 800
rect 344374 0 344430 800
rect 345478 0 345534 800
rect 346582 0 346638 800
rect 347686 0 347742 800
rect 348790 0 348846 800
rect 349894 0 349950 800
rect 350998 0 351054 800
rect 352102 0 352158 800
rect 353206 0 353262 800
rect 354310 0 354366 800
rect 355414 0 355470 800
rect 356518 0 356574 800
rect 357622 0 357678 800
rect 358726 0 358782 800
rect 359830 0 359886 800
rect 360934 0 360990 800
rect 362038 0 362094 800
rect 363142 0 363198 800
rect 364246 0 364302 800
rect 365350 0 365406 800
rect 366454 0 366510 800
rect 367558 0 367614 800
rect 368662 0 368718 800
rect 369766 0 369822 800
rect 370870 0 370926 800
rect 371974 0 372030 800
rect 373078 0 373134 800
rect 374182 0 374238 800
rect 375286 0 375342 800
rect 376390 0 376446 800
rect 377494 0 377550 800
rect 378598 0 378654 800
rect 379702 0 379758 800
rect 380806 0 380862 800
rect 381910 0 381966 800
rect 383014 0 383070 800
rect 384118 0 384174 800
rect 385222 0 385278 800
rect 386326 0 386382 800
rect 387430 0 387486 800
rect 388534 0 388590 800
rect 389638 0 389694 800
rect 390742 0 390798 800
rect 391846 0 391902 800
rect 392950 0 393006 800
rect 394054 0 394110 800
rect 395158 0 395214 800
rect 396262 0 396318 800
rect 397366 0 397422 800
rect 398470 0 398526 800
rect 399574 0 399630 800
rect 400678 0 400734 800
rect 401782 0 401838 800
rect 402886 0 402942 800
rect 403990 0 404046 800
rect 405094 0 405150 800
rect 406198 0 406254 800
rect 407302 0 407358 800
rect 408406 0 408462 800
rect 409510 0 409566 800
rect 410614 0 410670 800
rect 411718 0 411774 800
rect 412822 0 412878 800
rect 413926 0 413982 800
rect 415030 0 415086 800
rect 416134 0 416190 800
rect 417238 0 417294 800
rect 418342 0 418398 800
rect 419446 0 419502 800
rect 420550 0 420606 800
rect 421654 0 421710 800
rect 422758 0 422814 800
rect 423862 0 423918 800
rect 424966 0 425022 800
rect 426070 0 426126 800
rect 427174 0 427230 800
rect 428278 0 428334 800
rect 429382 0 429438 800
rect 430486 0 430542 800
rect 431590 0 431646 800
rect 432694 0 432750 800
rect 433798 0 433854 800
rect 434902 0 434958 800
rect 436006 0 436062 800
rect 437110 0 437166 800
rect 438214 0 438270 800
rect 439318 0 439374 800
rect 440422 0 440478 800
rect 441526 0 441582 800
rect 442630 0 442686 800
rect 443734 0 443790 800
rect 444838 0 444894 800
rect 445942 0 445998 800
rect 447046 0 447102 800
rect 448150 0 448206 800
rect 449254 0 449310 800
rect 450358 0 450414 800
rect 451462 0 451518 800
rect 452566 0 452622 800
rect 453670 0 453726 800
rect 454774 0 454830 800
rect 455878 0 455934 800
rect 456982 0 457038 800
rect 458086 0 458142 800
rect 459190 0 459246 800
rect 460294 0 460350 800
rect 461398 0 461454 800
rect 462502 0 462558 800
rect 463606 0 463662 800
rect 464710 0 464766 800
rect 465814 0 465870 800
rect 466918 0 466974 800
rect 468022 0 468078 800
rect 469126 0 469182 800
rect 470230 0 470286 800
rect 471334 0 471390 800
rect 472438 0 472494 800
rect 473542 0 473598 800
rect 474646 0 474702 800
rect 475750 0 475806 800
rect 476854 0 476910 800
rect 477958 0 478014 800
rect 479062 0 479118 800
rect 480166 0 480222 800
rect 481270 0 481326 800
rect 482374 0 482430 800
rect 483478 0 483534 800
rect 484582 0 484638 800
rect 485686 0 485742 800
rect 486790 0 486846 800
rect 487894 0 487950 800
rect 488998 0 489054 800
rect 490102 0 490158 800
rect 491206 0 491262 800
rect 492310 0 492366 800
rect 493414 0 493470 800
rect 494518 0 494574 800
rect 495622 0 495678 800
rect 496726 0 496782 800
rect 497830 0 497886 800
rect 498934 0 498990 800
rect 500038 0 500094 800
rect 501142 0 501198 800
rect 502246 0 502302 800
rect 503350 0 503406 800
rect 504454 0 504510 800
rect 505558 0 505614 800
rect 506662 0 506718 800
rect 507766 0 507822 800
rect 508870 0 508926 800
rect 509974 0 510030 800
rect 511078 0 511134 800
rect 512182 0 512238 800
rect 513286 0 513342 800
rect 514390 0 514446 800
rect 515494 0 515550 800
rect 516598 0 516654 800
rect 517702 0 517758 800
rect 518806 0 518862 800
rect 519910 0 519966 800
rect 521014 0 521070 800
rect 522118 0 522174 800
rect 523222 0 523278 800
rect 524326 0 524382 800
rect 525430 0 525486 800
rect 526534 0 526590 800
rect 527638 0 527694 800
rect 528742 0 528798 800
rect 529846 0 529902 800
rect 530950 0 531006 800
rect 532054 0 532110 800
rect 533158 0 533214 800
rect 534262 0 534318 800
rect 535366 0 535422 800
rect 536470 0 536526 800
rect 537574 0 537630 800
rect 538678 0 538734 800
rect 539782 0 539838 800
rect 540886 0 540942 800
rect 541990 0 542046 800
rect 543094 0 543150 800
rect 544198 0 544254 800
rect 545302 0 545358 800
rect 546406 0 546462 800
rect 547510 0 547566 800
rect 548614 0 548670 800
rect 549718 0 549774 800
rect 550822 0 550878 800
rect 551926 0 551982 800
rect 553030 0 553086 800
rect 554134 0 554190 800
rect 555238 0 555294 800
rect 556342 0 556398 800
rect 557446 0 557502 800
<< obsm2 >>
rect 386 685813 8334 685869
rect 8502 685813 24158 685869
rect 24326 685813 39982 685869
rect 40150 685813 55806 685869
rect 55974 685813 71630 685869
rect 71798 685813 87454 685869
rect 87622 685813 103278 685869
rect 103446 685813 119102 685869
rect 119270 685813 134926 685869
rect 135094 685813 150750 685869
rect 150918 685813 166574 685869
rect 166742 685813 182398 685869
rect 182566 685813 198222 685869
rect 198390 685813 214046 685869
rect 214214 685813 229870 685869
rect 230038 685813 245694 685869
rect 245862 685813 261518 685869
rect 261686 685813 277342 685869
rect 277510 685813 293166 685869
rect 293334 685813 308990 685869
rect 309158 685813 324814 685869
rect 324982 685813 340638 685869
rect 340806 685813 356462 685869
rect 356630 685813 372286 685869
rect 372454 685813 388110 685869
rect 388278 685813 403934 685869
rect 404102 685813 419758 685869
rect 419926 685813 435582 685869
rect 435750 685813 451406 685869
rect 451574 685813 467230 685869
rect 467398 685813 483054 685869
rect 483222 685813 498878 685869
rect 499046 685813 514702 685869
rect 514870 685813 530526 685869
rect 530694 685813 546350 685869
rect 546518 685813 562174 685869
rect 562342 685813 570748 685869
rect 386 856 570748 685813
rect 386 734 13118 856
rect 13286 734 14222 856
rect 14390 734 15326 856
rect 15494 734 16430 856
rect 16598 734 17534 856
rect 17702 734 18638 856
rect 18806 734 19742 856
rect 19910 734 20846 856
rect 21014 734 21950 856
rect 22118 734 23054 856
rect 23222 734 24158 856
rect 24326 734 25262 856
rect 25430 734 26366 856
rect 26534 734 27470 856
rect 27638 734 28574 856
rect 28742 734 29678 856
rect 29846 734 30782 856
rect 30950 734 31886 856
rect 32054 734 32990 856
rect 33158 734 34094 856
rect 34262 734 35198 856
rect 35366 734 36302 856
rect 36470 734 37406 856
rect 37574 734 38510 856
rect 38678 734 39614 856
rect 39782 734 40718 856
rect 40886 734 41822 856
rect 41990 734 42926 856
rect 43094 734 44030 856
rect 44198 734 45134 856
rect 45302 734 46238 856
rect 46406 734 47342 856
rect 47510 734 48446 856
rect 48614 734 49550 856
rect 49718 734 50654 856
rect 50822 734 51758 856
rect 51926 734 52862 856
rect 53030 734 53966 856
rect 54134 734 55070 856
rect 55238 734 56174 856
rect 56342 734 57278 856
rect 57446 734 58382 856
rect 58550 734 59486 856
rect 59654 734 60590 856
rect 60758 734 61694 856
rect 61862 734 62798 856
rect 62966 734 63902 856
rect 64070 734 65006 856
rect 65174 734 66110 856
rect 66278 734 67214 856
rect 67382 734 68318 856
rect 68486 734 69422 856
rect 69590 734 70526 856
rect 70694 734 71630 856
rect 71798 734 72734 856
rect 72902 734 73838 856
rect 74006 734 74942 856
rect 75110 734 76046 856
rect 76214 734 77150 856
rect 77318 734 78254 856
rect 78422 734 79358 856
rect 79526 734 80462 856
rect 80630 734 81566 856
rect 81734 734 82670 856
rect 82838 734 83774 856
rect 83942 734 84878 856
rect 85046 734 85982 856
rect 86150 734 87086 856
rect 87254 734 88190 856
rect 88358 734 89294 856
rect 89462 734 90398 856
rect 90566 734 91502 856
rect 91670 734 92606 856
rect 92774 734 93710 856
rect 93878 734 94814 856
rect 94982 734 95918 856
rect 96086 734 97022 856
rect 97190 734 98126 856
rect 98294 734 99230 856
rect 99398 734 100334 856
rect 100502 734 101438 856
rect 101606 734 102542 856
rect 102710 734 103646 856
rect 103814 734 104750 856
rect 104918 734 105854 856
rect 106022 734 106958 856
rect 107126 734 108062 856
rect 108230 734 109166 856
rect 109334 734 110270 856
rect 110438 734 111374 856
rect 111542 734 112478 856
rect 112646 734 113582 856
rect 113750 734 114686 856
rect 114854 734 115790 856
rect 115958 734 116894 856
rect 117062 734 117998 856
rect 118166 734 119102 856
rect 119270 734 120206 856
rect 120374 734 121310 856
rect 121478 734 122414 856
rect 122582 734 123518 856
rect 123686 734 124622 856
rect 124790 734 125726 856
rect 125894 734 126830 856
rect 126998 734 127934 856
rect 128102 734 129038 856
rect 129206 734 130142 856
rect 130310 734 131246 856
rect 131414 734 132350 856
rect 132518 734 133454 856
rect 133622 734 134558 856
rect 134726 734 135662 856
rect 135830 734 136766 856
rect 136934 734 137870 856
rect 138038 734 138974 856
rect 139142 734 140078 856
rect 140246 734 141182 856
rect 141350 734 142286 856
rect 142454 734 143390 856
rect 143558 734 144494 856
rect 144662 734 145598 856
rect 145766 734 146702 856
rect 146870 734 147806 856
rect 147974 734 148910 856
rect 149078 734 150014 856
rect 150182 734 151118 856
rect 151286 734 152222 856
rect 152390 734 153326 856
rect 153494 734 154430 856
rect 154598 734 155534 856
rect 155702 734 156638 856
rect 156806 734 157742 856
rect 157910 734 158846 856
rect 159014 734 159950 856
rect 160118 734 161054 856
rect 161222 734 162158 856
rect 162326 734 163262 856
rect 163430 734 164366 856
rect 164534 734 165470 856
rect 165638 734 166574 856
rect 166742 734 167678 856
rect 167846 734 168782 856
rect 168950 734 169886 856
rect 170054 734 170990 856
rect 171158 734 172094 856
rect 172262 734 173198 856
rect 173366 734 174302 856
rect 174470 734 175406 856
rect 175574 734 176510 856
rect 176678 734 177614 856
rect 177782 734 178718 856
rect 178886 734 179822 856
rect 179990 734 180926 856
rect 181094 734 182030 856
rect 182198 734 183134 856
rect 183302 734 184238 856
rect 184406 734 185342 856
rect 185510 734 186446 856
rect 186614 734 187550 856
rect 187718 734 188654 856
rect 188822 734 189758 856
rect 189926 734 190862 856
rect 191030 734 191966 856
rect 192134 734 193070 856
rect 193238 734 194174 856
rect 194342 734 195278 856
rect 195446 734 196382 856
rect 196550 734 197486 856
rect 197654 734 198590 856
rect 198758 734 199694 856
rect 199862 734 200798 856
rect 200966 734 201902 856
rect 202070 734 203006 856
rect 203174 734 204110 856
rect 204278 734 205214 856
rect 205382 734 206318 856
rect 206486 734 207422 856
rect 207590 734 208526 856
rect 208694 734 209630 856
rect 209798 734 210734 856
rect 210902 734 211838 856
rect 212006 734 212942 856
rect 213110 734 214046 856
rect 214214 734 215150 856
rect 215318 734 216254 856
rect 216422 734 217358 856
rect 217526 734 218462 856
rect 218630 734 219566 856
rect 219734 734 220670 856
rect 220838 734 221774 856
rect 221942 734 222878 856
rect 223046 734 223982 856
rect 224150 734 225086 856
rect 225254 734 226190 856
rect 226358 734 227294 856
rect 227462 734 228398 856
rect 228566 734 229502 856
rect 229670 734 230606 856
rect 230774 734 231710 856
rect 231878 734 232814 856
rect 232982 734 233918 856
rect 234086 734 235022 856
rect 235190 734 236126 856
rect 236294 734 237230 856
rect 237398 734 238334 856
rect 238502 734 239438 856
rect 239606 734 240542 856
rect 240710 734 241646 856
rect 241814 734 242750 856
rect 242918 734 243854 856
rect 244022 734 244958 856
rect 245126 734 246062 856
rect 246230 734 247166 856
rect 247334 734 248270 856
rect 248438 734 249374 856
rect 249542 734 250478 856
rect 250646 734 251582 856
rect 251750 734 252686 856
rect 252854 734 253790 856
rect 253958 734 254894 856
rect 255062 734 255998 856
rect 256166 734 257102 856
rect 257270 734 258206 856
rect 258374 734 259310 856
rect 259478 734 260414 856
rect 260582 734 261518 856
rect 261686 734 262622 856
rect 262790 734 263726 856
rect 263894 734 264830 856
rect 264998 734 265934 856
rect 266102 734 267038 856
rect 267206 734 268142 856
rect 268310 734 269246 856
rect 269414 734 270350 856
rect 270518 734 271454 856
rect 271622 734 272558 856
rect 272726 734 273662 856
rect 273830 734 274766 856
rect 274934 734 275870 856
rect 276038 734 276974 856
rect 277142 734 278078 856
rect 278246 734 279182 856
rect 279350 734 280286 856
rect 280454 734 281390 856
rect 281558 734 282494 856
rect 282662 734 283598 856
rect 283766 734 284702 856
rect 284870 734 285806 856
rect 285974 734 286910 856
rect 287078 734 288014 856
rect 288182 734 289118 856
rect 289286 734 290222 856
rect 290390 734 291326 856
rect 291494 734 292430 856
rect 292598 734 293534 856
rect 293702 734 294638 856
rect 294806 734 295742 856
rect 295910 734 296846 856
rect 297014 734 297950 856
rect 298118 734 299054 856
rect 299222 734 300158 856
rect 300326 734 301262 856
rect 301430 734 302366 856
rect 302534 734 303470 856
rect 303638 734 304574 856
rect 304742 734 305678 856
rect 305846 734 306782 856
rect 306950 734 307886 856
rect 308054 734 308990 856
rect 309158 734 310094 856
rect 310262 734 311198 856
rect 311366 734 312302 856
rect 312470 734 313406 856
rect 313574 734 314510 856
rect 314678 734 315614 856
rect 315782 734 316718 856
rect 316886 734 317822 856
rect 317990 734 318926 856
rect 319094 734 320030 856
rect 320198 734 321134 856
rect 321302 734 322238 856
rect 322406 734 323342 856
rect 323510 734 324446 856
rect 324614 734 325550 856
rect 325718 734 326654 856
rect 326822 734 327758 856
rect 327926 734 328862 856
rect 329030 734 329966 856
rect 330134 734 331070 856
rect 331238 734 332174 856
rect 332342 734 333278 856
rect 333446 734 334382 856
rect 334550 734 335486 856
rect 335654 734 336590 856
rect 336758 734 337694 856
rect 337862 734 338798 856
rect 338966 734 339902 856
rect 340070 734 341006 856
rect 341174 734 342110 856
rect 342278 734 343214 856
rect 343382 734 344318 856
rect 344486 734 345422 856
rect 345590 734 346526 856
rect 346694 734 347630 856
rect 347798 734 348734 856
rect 348902 734 349838 856
rect 350006 734 350942 856
rect 351110 734 352046 856
rect 352214 734 353150 856
rect 353318 734 354254 856
rect 354422 734 355358 856
rect 355526 734 356462 856
rect 356630 734 357566 856
rect 357734 734 358670 856
rect 358838 734 359774 856
rect 359942 734 360878 856
rect 361046 734 361982 856
rect 362150 734 363086 856
rect 363254 734 364190 856
rect 364358 734 365294 856
rect 365462 734 366398 856
rect 366566 734 367502 856
rect 367670 734 368606 856
rect 368774 734 369710 856
rect 369878 734 370814 856
rect 370982 734 371918 856
rect 372086 734 373022 856
rect 373190 734 374126 856
rect 374294 734 375230 856
rect 375398 734 376334 856
rect 376502 734 377438 856
rect 377606 734 378542 856
rect 378710 734 379646 856
rect 379814 734 380750 856
rect 380918 734 381854 856
rect 382022 734 382958 856
rect 383126 734 384062 856
rect 384230 734 385166 856
rect 385334 734 386270 856
rect 386438 734 387374 856
rect 387542 734 388478 856
rect 388646 734 389582 856
rect 389750 734 390686 856
rect 390854 734 391790 856
rect 391958 734 392894 856
rect 393062 734 393998 856
rect 394166 734 395102 856
rect 395270 734 396206 856
rect 396374 734 397310 856
rect 397478 734 398414 856
rect 398582 734 399518 856
rect 399686 734 400622 856
rect 400790 734 401726 856
rect 401894 734 402830 856
rect 402998 734 403934 856
rect 404102 734 405038 856
rect 405206 734 406142 856
rect 406310 734 407246 856
rect 407414 734 408350 856
rect 408518 734 409454 856
rect 409622 734 410558 856
rect 410726 734 411662 856
rect 411830 734 412766 856
rect 412934 734 413870 856
rect 414038 734 414974 856
rect 415142 734 416078 856
rect 416246 734 417182 856
rect 417350 734 418286 856
rect 418454 734 419390 856
rect 419558 734 420494 856
rect 420662 734 421598 856
rect 421766 734 422702 856
rect 422870 734 423806 856
rect 423974 734 424910 856
rect 425078 734 426014 856
rect 426182 734 427118 856
rect 427286 734 428222 856
rect 428390 734 429326 856
rect 429494 734 430430 856
rect 430598 734 431534 856
rect 431702 734 432638 856
rect 432806 734 433742 856
rect 433910 734 434846 856
rect 435014 734 435950 856
rect 436118 734 437054 856
rect 437222 734 438158 856
rect 438326 734 439262 856
rect 439430 734 440366 856
rect 440534 734 441470 856
rect 441638 734 442574 856
rect 442742 734 443678 856
rect 443846 734 444782 856
rect 444950 734 445886 856
rect 446054 734 446990 856
rect 447158 734 448094 856
rect 448262 734 449198 856
rect 449366 734 450302 856
rect 450470 734 451406 856
rect 451574 734 452510 856
rect 452678 734 453614 856
rect 453782 734 454718 856
rect 454886 734 455822 856
rect 455990 734 456926 856
rect 457094 734 458030 856
rect 458198 734 459134 856
rect 459302 734 460238 856
rect 460406 734 461342 856
rect 461510 734 462446 856
rect 462614 734 463550 856
rect 463718 734 464654 856
rect 464822 734 465758 856
rect 465926 734 466862 856
rect 467030 734 467966 856
rect 468134 734 469070 856
rect 469238 734 470174 856
rect 470342 734 471278 856
rect 471446 734 472382 856
rect 472550 734 473486 856
rect 473654 734 474590 856
rect 474758 734 475694 856
rect 475862 734 476798 856
rect 476966 734 477902 856
rect 478070 734 479006 856
rect 479174 734 480110 856
rect 480278 734 481214 856
rect 481382 734 482318 856
rect 482486 734 483422 856
rect 483590 734 484526 856
rect 484694 734 485630 856
rect 485798 734 486734 856
rect 486902 734 487838 856
rect 488006 734 488942 856
rect 489110 734 490046 856
rect 490214 734 491150 856
rect 491318 734 492254 856
rect 492422 734 493358 856
rect 493526 734 494462 856
rect 494630 734 495566 856
rect 495734 734 496670 856
rect 496838 734 497774 856
rect 497942 734 498878 856
rect 499046 734 499982 856
rect 500150 734 501086 856
rect 501254 734 502190 856
rect 502358 734 503294 856
rect 503462 734 504398 856
rect 504566 734 505502 856
rect 505670 734 506606 856
rect 506774 734 507710 856
rect 507878 734 508814 856
rect 508982 734 509918 856
rect 510086 734 511022 856
rect 511190 734 512126 856
rect 512294 734 513230 856
rect 513398 734 514334 856
rect 514502 734 515438 856
rect 515606 734 516542 856
rect 516710 734 517646 856
rect 517814 734 518750 856
rect 518918 734 519854 856
rect 520022 734 520958 856
rect 521126 734 522062 856
rect 522230 734 523166 856
rect 523334 734 524270 856
rect 524438 734 525374 856
rect 525542 734 526478 856
rect 526646 734 527582 856
rect 527750 734 528686 856
rect 528854 734 529790 856
rect 529958 734 530894 856
rect 531062 734 531998 856
rect 532166 734 533102 856
rect 533270 734 534206 856
rect 534374 734 535310 856
rect 535478 734 536414 856
rect 536582 734 537518 856
rect 537686 734 538622 856
rect 538790 734 539726 856
rect 539894 734 540830 856
rect 540998 734 541934 856
rect 542102 734 543038 856
rect 543206 734 544142 856
rect 544310 734 545246 856
rect 545414 734 546350 856
rect 546518 734 547454 856
rect 547622 734 548558 856
rect 548726 734 549662 856
rect 549830 734 550766 856
rect 550934 734 551870 856
rect 552038 734 552974 856
rect 553142 734 554078 856
rect 554246 734 555182 856
rect 555350 734 556286 856
rect 556454 734 557390 856
rect 557558 734 570748 856
<< metal3 >>
rect 570005 679192 570805 679312
rect 0 678376 800 678496
rect 570005 666272 570805 666392
rect 0 665728 800 665848
rect 570005 653352 570805 653472
rect 0 653080 800 653200
rect 0 640432 800 640552
rect 570005 640432 570805 640552
rect 0 627784 800 627904
rect 570005 627512 570805 627632
rect 0 615136 800 615256
rect 570005 614592 570805 614712
rect 0 602488 800 602608
rect 570005 601672 570805 601792
rect 0 589840 800 589960
rect 570005 588752 570805 588872
rect 0 577192 800 577312
rect 570005 575832 570805 575952
rect 0 564544 800 564664
rect 570005 562912 570805 563032
rect 0 551896 800 552016
rect 570005 549992 570805 550112
rect 0 539248 800 539368
rect 570005 537072 570805 537192
rect 0 526600 800 526720
rect 570005 524152 570805 524272
rect 0 513952 800 514072
rect 570005 511232 570805 511352
rect 0 501304 800 501424
rect 570005 498312 570805 498432
rect 0 488656 800 488776
rect 570005 485392 570805 485512
rect 0 476008 800 476128
rect 570005 472472 570805 472592
rect 0 463360 800 463480
rect 570005 459552 570805 459672
rect 0 450712 800 450832
rect 570005 446632 570805 446752
rect 0 438064 800 438184
rect 570005 433712 570805 433832
rect 0 425416 800 425536
rect 570005 420792 570805 420912
rect 0 412768 800 412888
rect 570005 407872 570805 407992
rect 0 400120 800 400240
rect 570005 394952 570805 395072
rect 0 387472 800 387592
rect 570005 382032 570805 382152
rect 0 374824 800 374944
rect 570005 369112 570805 369232
rect 0 362176 800 362296
rect 570005 356192 570805 356312
rect 0 349528 800 349648
rect 570005 343272 570805 343392
rect 0 336880 800 337000
rect 570005 330352 570805 330472
rect 0 324232 800 324352
rect 570005 317432 570805 317552
rect 0 311584 800 311704
rect 570005 304512 570805 304632
rect 0 298936 800 299056
rect 570005 291592 570805 291712
rect 0 286288 800 286408
rect 570005 278672 570805 278792
rect 0 273640 800 273760
rect 570005 265752 570805 265872
rect 0 260992 800 261112
rect 570005 252832 570805 252952
rect 0 248344 800 248464
rect 570005 239912 570805 240032
rect 0 235696 800 235816
rect 570005 226992 570805 227112
rect 0 223048 800 223168
rect 570005 214072 570805 214192
rect 0 210400 800 210520
rect 570005 201152 570805 201272
rect 0 197752 800 197872
rect 570005 188232 570805 188352
rect 0 185104 800 185224
rect 570005 175312 570805 175432
rect 0 172456 800 172576
rect 570005 162392 570805 162512
rect 0 159808 800 159928
rect 570005 149472 570805 149592
rect 0 147160 800 147280
rect 570005 136552 570805 136672
rect 0 134512 800 134632
rect 570005 123632 570805 123752
rect 0 121864 800 121984
rect 570005 110712 570805 110832
rect 0 109216 800 109336
rect 570005 97792 570805 97912
rect 0 96568 800 96688
rect 570005 84872 570805 84992
rect 0 83920 800 84040
rect 570005 71952 570805 72072
rect 0 71272 800 71392
rect 570005 59032 570805 59152
rect 0 58624 800 58744
rect 0 45976 800 46096
rect 570005 46112 570805 46232
rect 0 33328 800 33448
rect 570005 33192 570805 33312
rect 0 20680 800 20800
rect 570005 20272 570805 20392
rect 0 8032 800 8152
rect 570005 7352 570805 7472
<< obsm3 >>
rect 381 679392 570663 684385
rect 381 679112 569925 679392
rect 381 678576 570663 679112
rect 880 678296 570663 678576
rect 381 666472 570663 678296
rect 381 666192 569925 666472
rect 381 665928 570663 666192
rect 880 665648 570663 665928
rect 381 653552 570663 665648
rect 381 653280 569925 653552
rect 880 653272 569925 653280
rect 880 653000 570663 653272
rect 381 640632 570663 653000
rect 880 640352 569925 640632
rect 381 627984 570663 640352
rect 880 627712 570663 627984
rect 880 627704 569925 627712
rect 381 627432 569925 627704
rect 381 615336 570663 627432
rect 880 615056 570663 615336
rect 381 614792 570663 615056
rect 381 614512 569925 614792
rect 381 602688 570663 614512
rect 880 602408 570663 602688
rect 381 601872 570663 602408
rect 381 601592 569925 601872
rect 381 590040 570663 601592
rect 880 589760 570663 590040
rect 381 588952 570663 589760
rect 381 588672 569925 588952
rect 381 577392 570663 588672
rect 880 577112 570663 577392
rect 381 576032 570663 577112
rect 381 575752 569925 576032
rect 381 564744 570663 575752
rect 880 564464 570663 564744
rect 381 563112 570663 564464
rect 381 562832 569925 563112
rect 381 552096 570663 562832
rect 880 551816 570663 552096
rect 381 550192 570663 551816
rect 381 549912 569925 550192
rect 381 539448 570663 549912
rect 880 539168 570663 539448
rect 381 537272 570663 539168
rect 381 536992 569925 537272
rect 381 526800 570663 536992
rect 880 526520 570663 526800
rect 381 524352 570663 526520
rect 381 524072 569925 524352
rect 381 514152 570663 524072
rect 880 513872 570663 514152
rect 381 511432 570663 513872
rect 381 511152 569925 511432
rect 381 501504 570663 511152
rect 880 501224 570663 501504
rect 381 498512 570663 501224
rect 381 498232 569925 498512
rect 381 488856 570663 498232
rect 880 488576 570663 488856
rect 381 485592 570663 488576
rect 381 485312 569925 485592
rect 381 476208 570663 485312
rect 880 475928 570663 476208
rect 381 472672 570663 475928
rect 381 472392 569925 472672
rect 381 463560 570663 472392
rect 880 463280 570663 463560
rect 381 459752 570663 463280
rect 381 459472 569925 459752
rect 381 450912 570663 459472
rect 880 450632 570663 450912
rect 381 446832 570663 450632
rect 381 446552 569925 446832
rect 381 438264 570663 446552
rect 880 437984 570663 438264
rect 381 433912 570663 437984
rect 381 433632 569925 433912
rect 381 425616 570663 433632
rect 880 425336 570663 425616
rect 381 420992 570663 425336
rect 381 420712 569925 420992
rect 381 412968 570663 420712
rect 880 412688 570663 412968
rect 381 408072 570663 412688
rect 381 407792 569925 408072
rect 381 400320 570663 407792
rect 880 400040 570663 400320
rect 381 395152 570663 400040
rect 381 394872 569925 395152
rect 381 387672 570663 394872
rect 880 387392 570663 387672
rect 381 382232 570663 387392
rect 381 381952 569925 382232
rect 381 375024 570663 381952
rect 880 374744 570663 375024
rect 381 369312 570663 374744
rect 381 369032 569925 369312
rect 381 362376 570663 369032
rect 880 362096 570663 362376
rect 381 356392 570663 362096
rect 381 356112 569925 356392
rect 381 349728 570663 356112
rect 880 349448 570663 349728
rect 381 343472 570663 349448
rect 381 343192 569925 343472
rect 381 337080 570663 343192
rect 880 336800 570663 337080
rect 381 330552 570663 336800
rect 381 330272 569925 330552
rect 381 324432 570663 330272
rect 880 324152 570663 324432
rect 381 317632 570663 324152
rect 381 317352 569925 317632
rect 381 311784 570663 317352
rect 880 311504 570663 311784
rect 381 304712 570663 311504
rect 381 304432 569925 304712
rect 381 299136 570663 304432
rect 880 298856 570663 299136
rect 381 291792 570663 298856
rect 381 291512 569925 291792
rect 381 286488 570663 291512
rect 880 286208 570663 286488
rect 381 278872 570663 286208
rect 381 278592 569925 278872
rect 381 273840 570663 278592
rect 880 273560 570663 273840
rect 381 265952 570663 273560
rect 381 265672 569925 265952
rect 381 261192 570663 265672
rect 880 260912 570663 261192
rect 381 253032 570663 260912
rect 381 252752 569925 253032
rect 381 248544 570663 252752
rect 880 248264 570663 248544
rect 381 240112 570663 248264
rect 381 239832 569925 240112
rect 381 235896 570663 239832
rect 880 235616 570663 235896
rect 381 227192 570663 235616
rect 381 226912 569925 227192
rect 381 223248 570663 226912
rect 880 222968 570663 223248
rect 381 214272 570663 222968
rect 381 213992 569925 214272
rect 381 210600 570663 213992
rect 880 210320 570663 210600
rect 381 201352 570663 210320
rect 381 201072 569925 201352
rect 381 197952 570663 201072
rect 880 197672 570663 197952
rect 381 188432 570663 197672
rect 381 188152 569925 188432
rect 381 185304 570663 188152
rect 880 185024 570663 185304
rect 381 175512 570663 185024
rect 381 175232 569925 175512
rect 381 172656 570663 175232
rect 880 172376 570663 172656
rect 381 162592 570663 172376
rect 381 162312 569925 162592
rect 381 160008 570663 162312
rect 880 159728 570663 160008
rect 381 149672 570663 159728
rect 381 149392 569925 149672
rect 381 147360 570663 149392
rect 880 147080 570663 147360
rect 381 136752 570663 147080
rect 381 136472 569925 136752
rect 381 134712 570663 136472
rect 880 134432 570663 134712
rect 381 123832 570663 134432
rect 381 123552 569925 123832
rect 381 122064 570663 123552
rect 880 121784 570663 122064
rect 381 110912 570663 121784
rect 381 110632 569925 110912
rect 381 109416 570663 110632
rect 880 109136 570663 109416
rect 381 97992 570663 109136
rect 381 97712 569925 97992
rect 381 96768 570663 97712
rect 880 96488 570663 96768
rect 381 85072 570663 96488
rect 381 84792 569925 85072
rect 381 84120 570663 84792
rect 880 83840 570663 84120
rect 381 72152 570663 83840
rect 381 71872 569925 72152
rect 381 71472 570663 71872
rect 880 71192 570663 71472
rect 381 59232 570663 71192
rect 381 58952 569925 59232
rect 381 58824 570663 58952
rect 880 58544 570663 58824
rect 381 46312 570663 58544
rect 381 46176 569925 46312
rect 880 46032 569925 46176
rect 880 45896 570663 46032
rect 381 33528 570663 45896
rect 880 33392 570663 33528
rect 880 33248 569925 33392
rect 381 33112 569925 33248
rect 381 20880 570663 33112
rect 880 20600 570663 20880
rect 381 20472 570663 20600
rect 381 20192 569925 20472
rect 381 8232 570663 20192
rect 880 7952 570663 8232
rect 381 7552 570663 7952
rect 381 7272 569925 7552
rect 381 2143 570663 7272
<< metal4 >>
rect 4208 2128 4528 684400
rect 19568 2128 19888 684400
rect 34928 2128 35248 684400
rect 50288 2128 50608 684400
rect 65648 2128 65968 684400
rect 81008 2128 81328 684400
rect 96368 2128 96688 684400
rect 111728 2128 112048 684400
rect 127088 2128 127408 684400
rect 142448 2128 142768 684400
rect 157808 2128 158128 684400
rect 173168 2128 173488 684400
rect 188528 2128 188848 684400
rect 203888 2128 204208 684400
rect 219248 2128 219568 684400
rect 234608 2128 234928 684400
rect 249968 2128 250288 684400
rect 265328 2128 265648 684400
rect 280688 2128 281008 684400
rect 296048 2128 296368 684400
rect 311408 2128 311728 684400
rect 326768 2128 327088 684400
rect 342128 2128 342448 684400
rect 357488 2128 357808 684400
rect 372848 2128 373168 684400
rect 388208 2128 388528 684400
rect 403568 2128 403888 684400
rect 418928 2128 419248 684400
rect 434288 2128 434608 684400
rect 449648 2128 449968 684400
rect 465008 2128 465328 684400
rect 480368 2128 480688 684400
rect 495728 2128 496048 684400
rect 511088 2128 511408 684400
rect 526448 2128 526768 684400
rect 541808 2128 542128 684400
rect 557168 2128 557488 684400
<< obsm4 >>
rect 427 3435 4128 684045
rect 4608 3435 19488 684045
rect 19968 3435 34848 684045
rect 35328 3435 50208 684045
rect 50688 3435 65568 684045
rect 66048 3435 80928 684045
rect 81408 3435 96288 684045
rect 96768 3435 111648 684045
rect 112128 3435 127008 684045
rect 127488 3435 142368 684045
rect 142848 3435 157728 684045
rect 158208 3435 173088 684045
rect 173568 3435 188448 684045
rect 188928 3435 203808 684045
rect 204288 3435 219168 684045
rect 219648 3435 234528 684045
rect 235008 3435 249888 684045
rect 250368 3435 265248 684045
rect 265728 3435 280608 684045
rect 281088 3435 295968 684045
rect 296448 3435 311328 684045
rect 311808 3435 326688 684045
rect 327168 3435 342048 684045
rect 342528 3435 357408 684045
rect 357888 3435 372768 684045
rect 373248 3435 388128 684045
rect 388608 3435 403488 684045
rect 403968 3435 418848 684045
rect 419328 3435 434208 684045
rect 434688 3435 449568 684045
rect 450048 3435 464928 684045
rect 465408 3435 480288 684045
rect 480768 3435 495648 684045
rect 496128 3435 511008 684045
rect 511488 3435 526368 684045
rect 526848 3435 541728 684045
rect 542208 3435 557088 684045
rect 557568 3435 568501 684045
<< labels >>
rlabel metal3 s 570005 278672 570805 278792 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal2 s 435638 685869 435694 686669 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 372342 685869 372398 686669 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal2 s 309046 685869 309102 686669 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 245750 685869 245806 686669 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 182454 685869 182510 686669 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 119158 685869 119214 686669 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 55862 685869 55918 686669 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal3 s 0 678376 800 678496 6 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal3 s 0 627784 800 627904 6 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal3 s 0 577192 800 577312 6 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal3 s 570005 330352 570805 330472 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s 0 526600 800 526720 6 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal3 s 0 476008 800 476128 6 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s 0 425416 800 425536 6 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal3 s 0 374824 800 374944 6 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s 0 324232 800 324352 6 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal3 s 0 273640 800 273760 6 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s 0 223048 800 223168 6 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s 0 172456 800 172576 6 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s 0 121864 800 121984 6 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 570005 382032 570805 382152 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s 570005 433712 570805 433832 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal3 s 570005 485392 570805 485512 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal3 s 570005 537072 570805 537192 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal3 s 570005 588752 570805 588872 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal3 s 570005 640432 570805 640552 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal2 s 562230 685869 562286 686669 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal2 s 498934 685869 498990 686669 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal3 s 570005 7352 570805 7472 6 io_in[0]
port 30 nsew signal input
rlabel metal3 s 570005 446632 570805 446752 6 io_in[10]
port 31 nsew signal input
rlabel metal3 s 570005 498312 570805 498432 6 io_in[11]
port 32 nsew signal input
rlabel metal3 s 570005 549992 570805 550112 6 io_in[12]
port 33 nsew signal input
rlabel metal3 s 570005 601672 570805 601792 6 io_in[13]
port 34 nsew signal input
rlabel metal3 s 570005 653352 570805 653472 6 io_in[14]
port 35 nsew signal input
rlabel metal2 s 546406 685869 546462 686669 6 io_in[15]
port 36 nsew signal input
rlabel metal2 s 483110 685869 483166 686669 6 io_in[16]
port 37 nsew signal input
rlabel metal2 s 419814 685869 419870 686669 6 io_in[17]
port 38 nsew signal input
rlabel metal2 s 356518 685869 356574 686669 6 io_in[18]
port 39 nsew signal input
rlabel metal2 s 293222 685869 293278 686669 6 io_in[19]
port 40 nsew signal input
rlabel metal3 s 570005 46112 570805 46232 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 229926 685869 229982 686669 6 io_in[20]
port 42 nsew signal input
rlabel metal2 s 166630 685869 166686 686669 6 io_in[21]
port 43 nsew signal input
rlabel metal2 s 103334 685869 103390 686669 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 40038 685869 40094 686669 6 io_in[23]
port 45 nsew signal input
rlabel metal3 s 0 665728 800 665848 6 io_in[24]
port 46 nsew signal input
rlabel metal3 s 0 615136 800 615256 6 io_in[25]
port 47 nsew signal input
rlabel metal3 s 0 564544 800 564664 6 io_in[26]
port 48 nsew signal input
rlabel metal3 s 0 513952 800 514072 6 io_in[27]
port 49 nsew signal input
rlabel metal3 s 0 463360 800 463480 6 io_in[28]
port 50 nsew signal input
rlabel metal3 s 0 412768 800 412888 6 io_in[29]
port 51 nsew signal input
rlabel metal3 s 570005 84872 570805 84992 6 io_in[2]
port 52 nsew signal input
rlabel metal3 s 0 362176 800 362296 6 io_in[30]
port 53 nsew signal input
rlabel metal3 s 0 311584 800 311704 6 io_in[31]
port 54 nsew signal input
rlabel metal3 s 0 260992 800 261112 6 io_in[32]
port 55 nsew signal input
rlabel metal3 s 0 210400 800 210520 6 io_in[33]
port 56 nsew signal input
rlabel metal3 s 0 159808 800 159928 6 io_in[34]
port 57 nsew signal input
rlabel metal3 s 0 109216 800 109336 6 io_in[35]
port 58 nsew signal input
rlabel metal3 s 0 71272 800 71392 6 io_in[36]
port 59 nsew signal input
rlabel metal3 s 0 33328 800 33448 6 io_in[37]
port 60 nsew signal input
rlabel metal3 s 570005 123632 570805 123752 6 io_in[3]
port 61 nsew signal input
rlabel metal3 s 570005 162392 570805 162512 6 io_in[4]
port 62 nsew signal input
rlabel metal3 s 570005 201152 570805 201272 6 io_in[5]
port 63 nsew signal input
rlabel metal3 s 570005 239912 570805 240032 6 io_in[6]
port 64 nsew signal input
rlabel metal3 s 570005 291592 570805 291712 6 io_in[7]
port 65 nsew signal input
rlabel metal3 s 570005 343272 570805 343392 6 io_in[8]
port 66 nsew signal input
rlabel metal3 s 570005 394952 570805 395072 6 io_in[9]
port 67 nsew signal input
rlabel metal3 s 570005 33192 570805 33312 6 io_oeb[0]
port 68 nsew signal output
rlabel metal3 s 570005 472472 570805 472592 6 io_oeb[10]
port 69 nsew signal output
rlabel metal3 s 570005 524152 570805 524272 6 io_oeb[11]
port 70 nsew signal output
rlabel metal3 s 570005 575832 570805 575952 6 io_oeb[12]
port 71 nsew signal output
rlabel metal3 s 570005 627512 570805 627632 6 io_oeb[13]
port 72 nsew signal output
rlabel metal3 s 570005 679192 570805 679312 6 io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 514758 685869 514814 686669 6 io_oeb[15]
port 74 nsew signal output
rlabel metal2 s 451462 685869 451518 686669 6 io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 388166 685869 388222 686669 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 324870 685869 324926 686669 6 io_oeb[18]
port 77 nsew signal output
rlabel metal2 s 261574 685869 261630 686669 6 io_oeb[19]
port 78 nsew signal output
rlabel metal3 s 570005 71952 570805 72072 6 io_oeb[1]
port 79 nsew signal output
rlabel metal2 s 198278 685869 198334 686669 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 134982 685869 135038 686669 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 71686 685869 71742 686669 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 8390 685869 8446 686669 6 io_oeb[23]
port 83 nsew signal output
rlabel metal3 s 0 640432 800 640552 6 io_oeb[24]
port 84 nsew signal output
rlabel metal3 s 0 589840 800 589960 6 io_oeb[25]
port 85 nsew signal output
rlabel metal3 s 0 539248 800 539368 6 io_oeb[26]
port 86 nsew signal output
rlabel metal3 s 0 488656 800 488776 6 io_oeb[27]
port 87 nsew signal output
rlabel metal3 s 0 438064 800 438184 6 io_oeb[28]
port 88 nsew signal output
rlabel metal3 s 0 387472 800 387592 6 io_oeb[29]
port 89 nsew signal output
rlabel metal3 s 570005 110712 570805 110832 6 io_oeb[2]
port 90 nsew signal output
rlabel metal3 s 0 336880 800 337000 6 io_oeb[30]
port 91 nsew signal output
rlabel metal3 s 0 286288 800 286408 6 io_oeb[31]
port 92 nsew signal output
rlabel metal3 s 0 235696 800 235816 6 io_oeb[32]
port 93 nsew signal output
rlabel metal3 s 0 185104 800 185224 6 io_oeb[33]
port 94 nsew signal output
rlabel metal3 s 0 134512 800 134632 6 io_oeb[34]
port 95 nsew signal output
rlabel metal3 s 0 83920 800 84040 6 io_oeb[35]
port 96 nsew signal output
rlabel metal3 s 0 45976 800 46096 6 io_oeb[36]
port 97 nsew signal output
rlabel metal3 s 0 8032 800 8152 6 io_oeb[37]
port 98 nsew signal output
rlabel metal3 s 570005 149472 570805 149592 6 io_oeb[3]
port 99 nsew signal output
rlabel metal3 s 570005 188232 570805 188352 6 io_oeb[4]
port 100 nsew signal output
rlabel metal3 s 570005 226992 570805 227112 6 io_oeb[5]
port 101 nsew signal output
rlabel metal3 s 570005 265752 570805 265872 6 io_oeb[6]
port 102 nsew signal output
rlabel metal3 s 570005 317432 570805 317552 6 io_oeb[7]
port 103 nsew signal output
rlabel metal3 s 570005 369112 570805 369232 6 io_oeb[8]
port 104 nsew signal output
rlabel metal3 s 570005 420792 570805 420912 6 io_oeb[9]
port 105 nsew signal output
rlabel metal3 s 570005 20272 570805 20392 6 io_out[0]
port 106 nsew signal output
rlabel metal3 s 570005 459552 570805 459672 6 io_out[10]
port 107 nsew signal output
rlabel metal3 s 570005 511232 570805 511352 6 io_out[11]
port 108 nsew signal output
rlabel metal3 s 570005 562912 570805 563032 6 io_out[12]
port 109 nsew signal output
rlabel metal3 s 570005 614592 570805 614712 6 io_out[13]
port 110 nsew signal output
rlabel metal3 s 570005 666272 570805 666392 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 530582 685869 530638 686669 6 io_out[15]
port 112 nsew signal output
rlabel metal2 s 467286 685869 467342 686669 6 io_out[16]
port 113 nsew signal output
rlabel metal2 s 403990 685869 404046 686669 6 io_out[17]
port 114 nsew signal output
rlabel metal2 s 340694 685869 340750 686669 6 io_out[18]
port 115 nsew signal output
rlabel metal2 s 277398 685869 277454 686669 6 io_out[19]
port 116 nsew signal output
rlabel metal3 s 570005 59032 570805 59152 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 214102 685869 214158 686669 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 150806 685869 150862 686669 6 io_out[21]
port 119 nsew signal output
rlabel metal2 s 87510 685869 87566 686669 6 io_out[22]
port 120 nsew signal output
rlabel metal2 s 24214 685869 24270 686669 6 io_out[23]
port 121 nsew signal output
rlabel metal3 s 0 653080 800 653200 6 io_out[24]
port 122 nsew signal output
rlabel metal3 s 0 602488 800 602608 6 io_out[25]
port 123 nsew signal output
rlabel metal3 s 0 551896 800 552016 6 io_out[26]
port 124 nsew signal output
rlabel metal3 s 0 501304 800 501424 6 io_out[27]
port 125 nsew signal output
rlabel metal3 s 0 450712 800 450832 6 io_out[28]
port 126 nsew signal output
rlabel metal3 s 0 400120 800 400240 6 io_out[29]
port 127 nsew signal output
rlabel metal3 s 570005 97792 570805 97912 6 io_out[2]
port 128 nsew signal output
rlabel metal3 s 0 349528 800 349648 6 io_out[30]
port 129 nsew signal output
rlabel metal3 s 0 298936 800 299056 6 io_out[31]
port 130 nsew signal output
rlabel metal3 s 0 248344 800 248464 6 io_out[32]
port 131 nsew signal output
rlabel metal3 s 0 197752 800 197872 6 io_out[33]
port 132 nsew signal output
rlabel metal3 s 0 147160 800 147280 6 io_out[34]
port 133 nsew signal output
rlabel metal3 s 0 96568 800 96688 6 io_out[35]
port 134 nsew signal output
rlabel metal3 s 0 58624 800 58744 6 io_out[36]
port 135 nsew signal output
rlabel metal3 s 0 20680 800 20800 6 io_out[37]
port 136 nsew signal output
rlabel metal3 s 570005 136552 570805 136672 6 io_out[3]
port 137 nsew signal output
rlabel metal3 s 570005 175312 570805 175432 6 io_out[4]
port 138 nsew signal output
rlabel metal3 s 570005 214072 570805 214192 6 io_out[5]
port 139 nsew signal output
rlabel metal3 s 570005 252832 570805 252952 6 io_out[6]
port 140 nsew signal output
rlabel metal3 s 570005 304512 570805 304632 6 io_out[7]
port 141 nsew signal output
rlabel metal3 s 570005 356192 570805 356312 6 io_out[8]
port 142 nsew signal output
rlabel metal3 s 570005 407872 570805 407992 6 io_out[9]
port 143 nsew signal output
rlabel metal2 s 130198 0 130254 800 6 la_data_in[0]
port 144 nsew signal input
rlabel metal2 s 461398 0 461454 800 6 la_data_in[100]
port 145 nsew signal input
rlabel metal2 s 464710 0 464766 800 6 la_data_in[101]
port 146 nsew signal input
rlabel metal2 s 468022 0 468078 800 6 la_data_in[102]
port 147 nsew signal input
rlabel metal2 s 471334 0 471390 800 6 la_data_in[103]
port 148 nsew signal input
rlabel metal2 s 474646 0 474702 800 6 la_data_in[104]
port 149 nsew signal input
rlabel metal2 s 477958 0 478014 800 6 la_data_in[105]
port 150 nsew signal input
rlabel metal2 s 481270 0 481326 800 6 la_data_in[106]
port 151 nsew signal input
rlabel metal2 s 484582 0 484638 800 6 la_data_in[107]
port 152 nsew signal input
rlabel metal2 s 487894 0 487950 800 6 la_data_in[108]
port 153 nsew signal input
rlabel metal2 s 491206 0 491262 800 6 la_data_in[109]
port 154 nsew signal input
rlabel metal2 s 163318 0 163374 800 6 la_data_in[10]
port 155 nsew signal input
rlabel metal2 s 494518 0 494574 800 6 la_data_in[110]
port 156 nsew signal input
rlabel metal2 s 497830 0 497886 800 6 la_data_in[111]
port 157 nsew signal input
rlabel metal2 s 501142 0 501198 800 6 la_data_in[112]
port 158 nsew signal input
rlabel metal2 s 504454 0 504510 800 6 la_data_in[113]
port 159 nsew signal input
rlabel metal2 s 507766 0 507822 800 6 la_data_in[114]
port 160 nsew signal input
rlabel metal2 s 511078 0 511134 800 6 la_data_in[115]
port 161 nsew signal input
rlabel metal2 s 514390 0 514446 800 6 la_data_in[116]
port 162 nsew signal input
rlabel metal2 s 517702 0 517758 800 6 la_data_in[117]
port 163 nsew signal input
rlabel metal2 s 521014 0 521070 800 6 la_data_in[118]
port 164 nsew signal input
rlabel metal2 s 524326 0 524382 800 6 la_data_in[119]
port 165 nsew signal input
rlabel metal2 s 166630 0 166686 800 6 la_data_in[11]
port 166 nsew signal input
rlabel metal2 s 527638 0 527694 800 6 la_data_in[120]
port 167 nsew signal input
rlabel metal2 s 530950 0 531006 800 6 la_data_in[121]
port 168 nsew signal input
rlabel metal2 s 534262 0 534318 800 6 la_data_in[122]
port 169 nsew signal input
rlabel metal2 s 537574 0 537630 800 6 la_data_in[123]
port 170 nsew signal input
rlabel metal2 s 540886 0 540942 800 6 la_data_in[124]
port 171 nsew signal input
rlabel metal2 s 544198 0 544254 800 6 la_data_in[125]
port 172 nsew signal input
rlabel metal2 s 547510 0 547566 800 6 la_data_in[126]
port 173 nsew signal input
rlabel metal2 s 550822 0 550878 800 6 la_data_in[127]
port 174 nsew signal input
rlabel metal2 s 169942 0 169998 800 6 la_data_in[12]
port 175 nsew signal input
rlabel metal2 s 173254 0 173310 800 6 la_data_in[13]
port 176 nsew signal input
rlabel metal2 s 176566 0 176622 800 6 la_data_in[14]
port 177 nsew signal input
rlabel metal2 s 179878 0 179934 800 6 la_data_in[15]
port 178 nsew signal input
rlabel metal2 s 183190 0 183246 800 6 la_data_in[16]
port 179 nsew signal input
rlabel metal2 s 186502 0 186558 800 6 la_data_in[17]
port 180 nsew signal input
rlabel metal2 s 189814 0 189870 800 6 la_data_in[18]
port 181 nsew signal input
rlabel metal2 s 193126 0 193182 800 6 la_data_in[19]
port 182 nsew signal input
rlabel metal2 s 133510 0 133566 800 6 la_data_in[1]
port 183 nsew signal input
rlabel metal2 s 196438 0 196494 800 6 la_data_in[20]
port 184 nsew signal input
rlabel metal2 s 199750 0 199806 800 6 la_data_in[21]
port 185 nsew signal input
rlabel metal2 s 203062 0 203118 800 6 la_data_in[22]
port 186 nsew signal input
rlabel metal2 s 206374 0 206430 800 6 la_data_in[23]
port 187 nsew signal input
rlabel metal2 s 209686 0 209742 800 6 la_data_in[24]
port 188 nsew signal input
rlabel metal2 s 212998 0 213054 800 6 la_data_in[25]
port 189 nsew signal input
rlabel metal2 s 216310 0 216366 800 6 la_data_in[26]
port 190 nsew signal input
rlabel metal2 s 219622 0 219678 800 6 la_data_in[27]
port 191 nsew signal input
rlabel metal2 s 222934 0 222990 800 6 la_data_in[28]
port 192 nsew signal input
rlabel metal2 s 226246 0 226302 800 6 la_data_in[29]
port 193 nsew signal input
rlabel metal2 s 136822 0 136878 800 6 la_data_in[2]
port 194 nsew signal input
rlabel metal2 s 229558 0 229614 800 6 la_data_in[30]
port 195 nsew signal input
rlabel metal2 s 232870 0 232926 800 6 la_data_in[31]
port 196 nsew signal input
rlabel metal2 s 236182 0 236238 800 6 la_data_in[32]
port 197 nsew signal input
rlabel metal2 s 239494 0 239550 800 6 la_data_in[33]
port 198 nsew signal input
rlabel metal2 s 242806 0 242862 800 6 la_data_in[34]
port 199 nsew signal input
rlabel metal2 s 246118 0 246174 800 6 la_data_in[35]
port 200 nsew signal input
rlabel metal2 s 249430 0 249486 800 6 la_data_in[36]
port 201 nsew signal input
rlabel metal2 s 252742 0 252798 800 6 la_data_in[37]
port 202 nsew signal input
rlabel metal2 s 256054 0 256110 800 6 la_data_in[38]
port 203 nsew signal input
rlabel metal2 s 259366 0 259422 800 6 la_data_in[39]
port 204 nsew signal input
rlabel metal2 s 140134 0 140190 800 6 la_data_in[3]
port 205 nsew signal input
rlabel metal2 s 262678 0 262734 800 6 la_data_in[40]
port 206 nsew signal input
rlabel metal2 s 265990 0 266046 800 6 la_data_in[41]
port 207 nsew signal input
rlabel metal2 s 269302 0 269358 800 6 la_data_in[42]
port 208 nsew signal input
rlabel metal2 s 272614 0 272670 800 6 la_data_in[43]
port 209 nsew signal input
rlabel metal2 s 275926 0 275982 800 6 la_data_in[44]
port 210 nsew signal input
rlabel metal2 s 279238 0 279294 800 6 la_data_in[45]
port 211 nsew signal input
rlabel metal2 s 282550 0 282606 800 6 la_data_in[46]
port 212 nsew signal input
rlabel metal2 s 285862 0 285918 800 6 la_data_in[47]
port 213 nsew signal input
rlabel metal2 s 289174 0 289230 800 6 la_data_in[48]
port 214 nsew signal input
rlabel metal2 s 292486 0 292542 800 6 la_data_in[49]
port 215 nsew signal input
rlabel metal2 s 143446 0 143502 800 6 la_data_in[4]
port 216 nsew signal input
rlabel metal2 s 295798 0 295854 800 6 la_data_in[50]
port 217 nsew signal input
rlabel metal2 s 299110 0 299166 800 6 la_data_in[51]
port 218 nsew signal input
rlabel metal2 s 302422 0 302478 800 6 la_data_in[52]
port 219 nsew signal input
rlabel metal2 s 305734 0 305790 800 6 la_data_in[53]
port 220 nsew signal input
rlabel metal2 s 309046 0 309102 800 6 la_data_in[54]
port 221 nsew signal input
rlabel metal2 s 312358 0 312414 800 6 la_data_in[55]
port 222 nsew signal input
rlabel metal2 s 315670 0 315726 800 6 la_data_in[56]
port 223 nsew signal input
rlabel metal2 s 318982 0 319038 800 6 la_data_in[57]
port 224 nsew signal input
rlabel metal2 s 322294 0 322350 800 6 la_data_in[58]
port 225 nsew signal input
rlabel metal2 s 325606 0 325662 800 6 la_data_in[59]
port 226 nsew signal input
rlabel metal2 s 146758 0 146814 800 6 la_data_in[5]
port 227 nsew signal input
rlabel metal2 s 328918 0 328974 800 6 la_data_in[60]
port 228 nsew signal input
rlabel metal2 s 332230 0 332286 800 6 la_data_in[61]
port 229 nsew signal input
rlabel metal2 s 335542 0 335598 800 6 la_data_in[62]
port 230 nsew signal input
rlabel metal2 s 338854 0 338910 800 6 la_data_in[63]
port 231 nsew signal input
rlabel metal2 s 342166 0 342222 800 6 la_data_in[64]
port 232 nsew signal input
rlabel metal2 s 345478 0 345534 800 6 la_data_in[65]
port 233 nsew signal input
rlabel metal2 s 348790 0 348846 800 6 la_data_in[66]
port 234 nsew signal input
rlabel metal2 s 352102 0 352158 800 6 la_data_in[67]
port 235 nsew signal input
rlabel metal2 s 355414 0 355470 800 6 la_data_in[68]
port 236 nsew signal input
rlabel metal2 s 358726 0 358782 800 6 la_data_in[69]
port 237 nsew signal input
rlabel metal2 s 150070 0 150126 800 6 la_data_in[6]
port 238 nsew signal input
rlabel metal2 s 362038 0 362094 800 6 la_data_in[70]
port 239 nsew signal input
rlabel metal2 s 365350 0 365406 800 6 la_data_in[71]
port 240 nsew signal input
rlabel metal2 s 368662 0 368718 800 6 la_data_in[72]
port 241 nsew signal input
rlabel metal2 s 371974 0 372030 800 6 la_data_in[73]
port 242 nsew signal input
rlabel metal2 s 375286 0 375342 800 6 la_data_in[74]
port 243 nsew signal input
rlabel metal2 s 378598 0 378654 800 6 la_data_in[75]
port 244 nsew signal input
rlabel metal2 s 381910 0 381966 800 6 la_data_in[76]
port 245 nsew signal input
rlabel metal2 s 385222 0 385278 800 6 la_data_in[77]
port 246 nsew signal input
rlabel metal2 s 388534 0 388590 800 6 la_data_in[78]
port 247 nsew signal input
rlabel metal2 s 391846 0 391902 800 6 la_data_in[79]
port 248 nsew signal input
rlabel metal2 s 153382 0 153438 800 6 la_data_in[7]
port 249 nsew signal input
rlabel metal2 s 395158 0 395214 800 6 la_data_in[80]
port 250 nsew signal input
rlabel metal2 s 398470 0 398526 800 6 la_data_in[81]
port 251 nsew signal input
rlabel metal2 s 401782 0 401838 800 6 la_data_in[82]
port 252 nsew signal input
rlabel metal2 s 405094 0 405150 800 6 la_data_in[83]
port 253 nsew signal input
rlabel metal2 s 408406 0 408462 800 6 la_data_in[84]
port 254 nsew signal input
rlabel metal2 s 411718 0 411774 800 6 la_data_in[85]
port 255 nsew signal input
rlabel metal2 s 415030 0 415086 800 6 la_data_in[86]
port 256 nsew signal input
rlabel metal2 s 418342 0 418398 800 6 la_data_in[87]
port 257 nsew signal input
rlabel metal2 s 421654 0 421710 800 6 la_data_in[88]
port 258 nsew signal input
rlabel metal2 s 424966 0 425022 800 6 la_data_in[89]
port 259 nsew signal input
rlabel metal2 s 156694 0 156750 800 6 la_data_in[8]
port 260 nsew signal input
rlabel metal2 s 428278 0 428334 800 6 la_data_in[90]
port 261 nsew signal input
rlabel metal2 s 431590 0 431646 800 6 la_data_in[91]
port 262 nsew signal input
rlabel metal2 s 434902 0 434958 800 6 la_data_in[92]
port 263 nsew signal input
rlabel metal2 s 438214 0 438270 800 6 la_data_in[93]
port 264 nsew signal input
rlabel metal2 s 441526 0 441582 800 6 la_data_in[94]
port 265 nsew signal input
rlabel metal2 s 444838 0 444894 800 6 la_data_in[95]
port 266 nsew signal input
rlabel metal2 s 448150 0 448206 800 6 la_data_in[96]
port 267 nsew signal input
rlabel metal2 s 451462 0 451518 800 6 la_data_in[97]
port 268 nsew signal input
rlabel metal2 s 454774 0 454830 800 6 la_data_in[98]
port 269 nsew signal input
rlabel metal2 s 458086 0 458142 800 6 la_data_in[99]
port 270 nsew signal input
rlabel metal2 s 160006 0 160062 800 6 la_data_in[9]
port 271 nsew signal input
rlabel metal2 s 131302 0 131358 800 6 la_data_out[0]
port 272 nsew signal output
rlabel metal2 s 462502 0 462558 800 6 la_data_out[100]
port 273 nsew signal output
rlabel metal2 s 465814 0 465870 800 6 la_data_out[101]
port 274 nsew signal output
rlabel metal2 s 469126 0 469182 800 6 la_data_out[102]
port 275 nsew signal output
rlabel metal2 s 472438 0 472494 800 6 la_data_out[103]
port 276 nsew signal output
rlabel metal2 s 475750 0 475806 800 6 la_data_out[104]
port 277 nsew signal output
rlabel metal2 s 479062 0 479118 800 6 la_data_out[105]
port 278 nsew signal output
rlabel metal2 s 482374 0 482430 800 6 la_data_out[106]
port 279 nsew signal output
rlabel metal2 s 485686 0 485742 800 6 la_data_out[107]
port 280 nsew signal output
rlabel metal2 s 488998 0 489054 800 6 la_data_out[108]
port 281 nsew signal output
rlabel metal2 s 492310 0 492366 800 6 la_data_out[109]
port 282 nsew signal output
rlabel metal2 s 164422 0 164478 800 6 la_data_out[10]
port 283 nsew signal output
rlabel metal2 s 495622 0 495678 800 6 la_data_out[110]
port 284 nsew signal output
rlabel metal2 s 498934 0 498990 800 6 la_data_out[111]
port 285 nsew signal output
rlabel metal2 s 502246 0 502302 800 6 la_data_out[112]
port 286 nsew signal output
rlabel metal2 s 505558 0 505614 800 6 la_data_out[113]
port 287 nsew signal output
rlabel metal2 s 508870 0 508926 800 6 la_data_out[114]
port 288 nsew signal output
rlabel metal2 s 512182 0 512238 800 6 la_data_out[115]
port 289 nsew signal output
rlabel metal2 s 515494 0 515550 800 6 la_data_out[116]
port 290 nsew signal output
rlabel metal2 s 518806 0 518862 800 6 la_data_out[117]
port 291 nsew signal output
rlabel metal2 s 522118 0 522174 800 6 la_data_out[118]
port 292 nsew signal output
rlabel metal2 s 525430 0 525486 800 6 la_data_out[119]
port 293 nsew signal output
rlabel metal2 s 167734 0 167790 800 6 la_data_out[11]
port 294 nsew signal output
rlabel metal2 s 528742 0 528798 800 6 la_data_out[120]
port 295 nsew signal output
rlabel metal2 s 532054 0 532110 800 6 la_data_out[121]
port 296 nsew signal output
rlabel metal2 s 535366 0 535422 800 6 la_data_out[122]
port 297 nsew signal output
rlabel metal2 s 538678 0 538734 800 6 la_data_out[123]
port 298 nsew signal output
rlabel metal2 s 541990 0 542046 800 6 la_data_out[124]
port 299 nsew signal output
rlabel metal2 s 545302 0 545358 800 6 la_data_out[125]
port 300 nsew signal output
rlabel metal2 s 548614 0 548670 800 6 la_data_out[126]
port 301 nsew signal output
rlabel metal2 s 551926 0 551982 800 6 la_data_out[127]
port 302 nsew signal output
rlabel metal2 s 171046 0 171102 800 6 la_data_out[12]
port 303 nsew signal output
rlabel metal2 s 174358 0 174414 800 6 la_data_out[13]
port 304 nsew signal output
rlabel metal2 s 177670 0 177726 800 6 la_data_out[14]
port 305 nsew signal output
rlabel metal2 s 180982 0 181038 800 6 la_data_out[15]
port 306 nsew signal output
rlabel metal2 s 184294 0 184350 800 6 la_data_out[16]
port 307 nsew signal output
rlabel metal2 s 187606 0 187662 800 6 la_data_out[17]
port 308 nsew signal output
rlabel metal2 s 190918 0 190974 800 6 la_data_out[18]
port 309 nsew signal output
rlabel metal2 s 194230 0 194286 800 6 la_data_out[19]
port 310 nsew signal output
rlabel metal2 s 134614 0 134670 800 6 la_data_out[1]
port 311 nsew signal output
rlabel metal2 s 197542 0 197598 800 6 la_data_out[20]
port 312 nsew signal output
rlabel metal2 s 200854 0 200910 800 6 la_data_out[21]
port 313 nsew signal output
rlabel metal2 s 204166 0 204222 800 6 la_data_out[22]
port 314 nsew signal output
rlabel metal2 s 207478 0 207534 800 6 la_data_out[23]
port 315 nsew signal output
rlabel metal2 s 210790 0 210846 800 6 la_data_out[24]
port 316 nsew signal output
rlabel metal2 s 214102 0 214158 800 6 la_data_out[25]
port 317 nsew signal output
rlabel metal2 s 217414 0 217470 800 6 la_data_out[26]
port 318 nsew signal output
rlabel metal2 s 220726 0 220782 800 6 la_data_out[27]
port 319 nsew signal output
rlabel metal2 s 224038 0 224094 800 6 la_data_out[28]
port 320 nsew signal output
rlabel metal2 s 227350 0 227406 800 6 la_data_out[29]
port 321 nsew signal output
rlabel metal2 s 137926 0 137982 800 6 la_data_out[2]
port 322 nsew signal output
rlabel metal2 s 230662 0 230718 800 6 la_data_out[30]
port 323 nsew signal output
rlabel metal2 s 233974 0 234030 800 6 la_data_out[31]
port 324 nsew signal output
rlabel metal2 s 237286 0 237342 800 6 la_data_out[32]
port 325 nsew signal output
rlabel metal2 s 240598 0 240654 800 6 la_data_out[33]
port 326 nsew signal output
rlabel metal2 s 243910 0 243966 800 6 la_data_out[34]
port 327 nsew signal output
rlabel metal2 s 247222 0 247278 800 6 la_data_out[35]
port 328 nsew signal output
rlabel metal2 s 250534 0 250590 800 6 la_data_out[36]
port 329 nsew signal output
rlabel metal2 s 253846 0 253902 800 6 la_data_out[37]
port 330 nsew signal output
rlabel metal2 s 257158 0 257214 800 6 la_data_out[38]
port 331 nsew signal output
rlabel metal2 s 260470 0 260526 800 6 la_data_out[39]
port 332 nsew signal output
rlabel metal2 s 141238 0 141294 800 6 la_data_out[3]
port 333 nsew signal output
rlabel metal2 s 263782 0 263838 800 6 la_data_out[40]
port 334 nsew signal output
rlabel metal2 s 267094 0 267150 800 6 la_data_out[41]
port 335 nsew signal output
rlabel metal2 s 270406 0 270462 800 6 la_data_out[42]
port 336 nsew signal output
rlabel metal2 s 273718 0 273774 800 6 la_data_out[43]
port 337 nsew signal output
rlabel metal2 s 277030 0 277086 800 6 la_data_out[44]
port 338 nsew signal output
rlabel metal2 s 280342 0 280398 800 6 la_data_out[45]
port 339 nsew signal output
rlabel metal2 s 283654 0 283710 800 6 la_data_out[46]
port 340 nsew signal output
rlabel metal2 s 286966 0 287022 800 6 la_data_out[47]
port 341 nsew signal output
rlabel metal2 s 290278 0 290334 800 6 la_data_out[48]
port 342 nsew signal output
rlabel metal2 s 293590 0 293646 800 6 la_data_out[49]
port 343 nsew signal output
rlabel metal2 s 144550 0 144606 800 6 la_data_out[4]
port 344 nsew signal output
rlabel metal2 s 296902 0 296958 800 6 la_data_out[50]
port 345 nsew signal output
rlabel metal2 s 300214 0 300270 800 6 la_data_out[51]
port 346 nsew signal output
rlabel metal2 s 303526 0 303582 800 6 la_data_out[52]
port 347 nsew signal output
rlabel metal2 s 306838 0 306894 800 6 la_data_out[53]
port 348 nsew signal output
rlabel metal2 s 310150 0 310206 800 6 la_data_out[54]
port 349 nsew signal output
rlabel metal2 s 313462 0 313518 800 6 la_data_out[55]
port 350 nsew signal output
rlabel metal2 s 316774 0 316830 800 6 la_data_out[56]
port 351 nsew signal output
rlabel metal2 s 320086 0 320142 800 6 la_data_out[57]
port 352 nsew signal output
rlabel metal2 s 323398 0 323454 800 6 la_data_out[58]
port 353 nsew signal output
rlabel metal2 s 326710 0 326766 800 6 la_data_out[59]
port 354 nsew signal output
rlabel metal2 s 147862 0 147918 800 6 la_data_out[5]
port 355 nsew signal output
rlabel metal2 s 330022 0 330078 800 6 la_data_out[60]
port 356 nsew signal output
rlabel metal2 s 333334 0 333390 800 6 la_data_out[61]
port 357 nsew signal output
rlabel metal2 s 336646 0 336702 800 6 la_data_out[62]
port 358 nsew signal output
rlabel metal2 s 339958 0 340014 800 6 la_data_out[63]
port 359 nsew signal output
rlabel metal2 s 343270 0 343326 800 6 la_data_out[64]
port 360 nsew signal output
rlabel metal2 s 346582 0 346638 800 6 la_data_out[65]
port 361 nsew signal output
rlabel metal2 s 349894 0 349950 800 6 la_data_out[66]
port 362 nsew signal output
rlabel metal2 s 353206 0 353262 800 6 la_data_out[67]
port 363 nsew signal output
rlabel metal2 s 356518 0 356574 800 6 la_data_out[68]
port 364 nsew signal output
rlabel metal2 s 359830 0 359886 800 6 la_data_out[69]
port 365 nsew signal output
rlabel metal2 s 151174 0 151230 800 6 la_data_out[6]
port 366 nsew signal output
rlabel metal2 s 363142 0 363198 800 6 la_data_out[70]
port 367 nsew signal output
rlabel metal2 s 366454 0 366510 800 6 la_data_out[71]
port 368 nsew signal output
rlabel metal2 s 369766 0 369822 800 6 la_data_out[72]
port 369 nsew signal output
rlabel metal2 s 373078 0 373134 800 6 la_data_out[73]
port 370 nsew signal output
rlabel metal2 s 376390 0 376446 800 6 la_data_out[74]
port 371 nsew signal output
rlabel metal2 s 379702 0 379758 800 6 la_data_out[75]
port 372 nsew signal output
rlabel metal2 s 383014 0 383070 800 6 la_data_out[76]
port 373 nsew signal output
rlabel metal2 s 386326 0 386382 800 6 la_data_out[77]
port 374 nsew signal output
rlabel metal2 s 389638 0 389694 800 6 la_data_out[78]
port 375 nsew signal output
rlabel metal2 s 392950 0 393006 800 6 la_data_out[79]
port 376 nsew signal output
rlabel metal2 s 154486 0 154542 800 6 la_data_out[7]
port 377 nsew signal output
rlabel metal2 s 396262 0 396318 800 6 la_data_out[80]
port 378 nsew signal output
rlabel metal2 s 399574 0 399630 800 6 la_data_out[81]
port 379 nsew signal output
rlabel metal2 s 402886 0 402942 800 6 la_data_out[82]
port 380 nsew signal output
rlabel metal2 s 406198 0 406254 800 6 la_data_out[83]
port 381 nsew signal output
rlabel metal2 s 409510 0 409566 800 6 la_data_out[84]
port 382 nsew signal output
rlabel metal2 s 412822 0 412878 800 6 la_data_out[85]
port 383 nsew signal output
rlabel metal2 s 416134 0 416190 800 6 la_data_out[86]
port 384 nsew signal output
rlabel metal2 s 419446 0 419502 800 6 la_data_out[87]
port 385 nsew signal output
rlabel metal2 s 422758 0 422814 800 6 la_data_out[88]
port 386 nsew signal output
rlabel metal2 s 426070 0 426126 800 6 la_data_out[89]
port 387 nsew signal output
rlabel metal2 s 157798 0 157854 800 6 la_data_out[8]
port 388 nsew signal output
rlabel metal2 s 429382 0 429438 800 6 la_data_out[90]
port 389 nsew signal output
rlabel metal2 s 432694 0 432750 800 6 la_data_out[91]
port 390 nsew signal output
rlabel metal2 s 436006 0 436062 800 6 la_data_out[92]
port 391 nsew signal output
rlabel metal2 s 439318 0 439374 800 6 la_data_out[93]
port 392 nsew signal output
rlabel metal2 s 442630 0 442686 800 6 la_data_out[94]
port 393 nsew signal output
rlabel metal2 s 445942 0 445998 800 6 la_data_out[95]
port 394 nsew signal output
rlabel metal2 s 449254 0 449310 800 6 la_data_out[96]
port 395 nsew signal output
rlabel metal2 s 452566 0 452622 800 6 la_data_out[97]
port 396 nsew signal output
rlabel metal2 s 455878 0 455934 800 6 la_data_out[98]
port 397 nsew signal output
rlabel metal2 s 459190 0 459246 800 6 la_data_out[99]
port 398 nsew signal output
rlabel metal2 s 161110 0 161166 800 6 la_data_out[9]
port 399 nsew signal output
rlabel metal2 s 132406 0 132462 800 6 la_oenb[0]
port 400 nsew signal input
rlabel metal2 s 463606 0 463662 800 6 la_oenb[100]
port 401 nsew signal input
rlabel metal2 s 466918 0 466974 800 6 la_oenb[101]
port 402 nsew signal input
rlabel metal2 s 470230 0 470286 800 6 la_oenb[102]
port 403 nsew signal input
rlabel metal2 s 473542 0 473598 800 6 la_oenb[103]
port 404 nsew signal input
rlabel metal2 s 476854 0 476910 800 6 la_oenb[104]
port 405 nsew signal input
rlabel metal2 s 480166 0 480222 800 6 la_oenb[105]
port 406 nsew signal input
rlabel metal2 s 483478 0 483534 800 6 la_oenb[106]
port 407 nsew signal input
rlabel metal2 s 486790 0 486846 800 6 la_oenb[107]
port 408 nsew signal input
rlabel metal2 s 490102 0 490158 800 6 la_oenb[108]
port 409 nsew signal input
rlabel metal2 s 493414 0 493470 800 6 la_oenb[109]
port 410 nsew signal input
rlabel metal2 s 165526 0 165582 800 6 la_oenb[10]
port 411 nsew signal input
rlabel metal2 s 496726 0 496782 800 6 la_oenb[110]
port 412 nsew signal input
rlabel metal2 s 500038 0 500094 800 6 la_oenb[111]
port 413 nsew signal input
rlabel metal2 s 503350 0 503406 800 6 la_oenb[112]
port 414 nsew signal input
rlabel metal2 s 506662 0 506718 800 6 la_oenb[113]
port 415 nsew signal input
rlabel metal2 s 509974 0 510030 800 6 la_oenb[114]
port 416 nsew signal input
rlabel metal2 s 513286 0 513342 800 6 la_oenb[115]
port 417 nsew signal input
rlabel metal2 s 516598 0 516654 800 6 la_oenb[116]
port 418 nsew signal input
rlabel metal2 s 519910 0 519966 800 6 la_oenb[117]
port 419 nsew signal input
rlabel metal2 s 523222 0 523278 800 6 la_oenb[118]
port 420 nsew signal input
rlabel metal2 s 526534 0 526590 800 6 la_oenb[119]
port 421 nsew signal input
rlabel metal2 s 168838 0 168894 800 6 la_oenb[11]
port 422 nsew signal input
rlabel metal2 s 529846 0 529902 800 6 la_oenb[120]
port 423 nsew signal input
rlabel metal2 s 533158 0 533214 800 6 la_oenb[121]
port 424 nsew signal input
rlabel metal2 s 536470 0 536526 800 6 la_oenb[122]
port 425 nsew signal input
rlabel metal2 s 539782 0 539838 800 6 la_oenb[123]
port 426 nsew signal input
rlabel metal2 s 543094 0 543150 800 6 la_oenb[124]
port 427 nsew signal input
rlabel metal2 s 546406 0 546462 800 6 la_oenb[125]
port 428 nsew signal input
rlabel metal2 s 549718 0 549774 800 6 la_oenb[126]
port 429 nsew signal input
rlabel metal2 s 553030 0 553086 800 6 la_oenb[127]
port 430 nsew signal input
rlabel metal2 s 172150 0 172206 800 6 la_oenb[12]
port 431 nsew signal input
rlabel metal2 s 175462 0 175518 800 6 la_oenb[13]
port 432 nsew signal input
rlabel metal2 s 178774 0 178830 800 6 la_oenb[14]
port 433 nsew signal input
rlabel metal2 s 182086 0 182142 800 6 la_oenb[15]
port 434 nsew signal input
rlabel metal2 s 185398 0 185454 800 6 la_oenb[16]
port 435 nsew signal input
rlabel metal2 s 188710 0 188766 800 6 la_oenb[17]
port 436 nsew signal input
rlabel metal2 s 192022 0 192078 800 6 la_oenb[18]
port 437 nsew signal input
rlabel metal2 s 195334 0 195390 800 6 la_oenb[19]
port 438 nsew signal input
rlabel metal2 s 135718 0 135774 800 6 la_oenb[1]
port 439 nsew signal input
rlabel metal2 s 198646 0 198702 800 6 la_oenb[20]
port 440 nsew signal input
rlabel metal2 s 201958 0 202014 800 6 la_oenb[21]
port 441 nsew signal input
rlabel metal2 s 205270 0 205326 800 6 la_oenb[22]
port 442 nsew signal input
rlabel metal2 s 208582 0 208638 800 6 la_oenb[23]
port 443 nsew signal input
rlabel metal2 s 211894 0 211950 800 6 la_oenb[24]
port 444 nsew signal input
rlabel metal2 s 215206 0 215262 800 6 la_oenb[25]
port 445 nsew signal input
rlabel metal2 s 218518 0 218574 800 6 la_oenb[26]
port 446 nsew signal input
rlabel metal2 s 221830 0 221886 800 6 la_oenb[27]
port 447 nsew signal input
rlabel metal2 s 225142 0 225198 800 6 la_oenb[28]
port 448 nsew signal input
rlabel metal2 s 228454 0 228510 800 6 la_oenb[29]
port 449 nsew signal input
rlabel metal2 s 139030 0 139086 800 6 la_oenb[2]
port 450 nsew signal input
rlabel metal2 s 231766 0 231822 800 6 la_oenb[30]
port 451 nsew signal input
rlabel metal2 s 235078 0 235134 800 6 la_oenb[31]
port 452 nsew signal input
rlabel metal2 s 238390 0 238446 800 6 la_oenb[32]
port 453 nsew signal input
rlabel metal2 s 241702 0 241758 800 6 la_oenb[33]
port 454 nsew signal input
rlabel metal2 s 245014 0 245070 800 6 la_oenb[34]
port 455 nsew signal input
rlabel metal2 s 248326 0 248382 800 6 la_oenb[35]
port 456 nsew signal input
rlabel metal2 s 251638 0 251694 800 6 la_oenb[36]
port 457 nsew signal input
rlabel metal2 s 254950 0 255006 800 6 la_oenb[37]
port 458 nsew signal input
rlabel metal2 s 258262 0 258318 800 6 la_oenb[38]
port 459 nsew signal input
rlabel metal2 s 261574 0 261630 800 6 la_oenb[39]
port 460 nsew signal input
rlabel metal2 s 142342 0 142398 800 6 la_oenb[3]
port 461 nsew signal input
rlabel metal2 s 264886 0 264942 800 6 la_oenb[40]
port 462 nsew signal input
rlabel metal2 s 268198 0 268254 800 6 la_oenb[41]
port 463 nsew signal input
rlabel metal2 s 271510 0 271566 800 6 la_oenb[42]
port 464 nsew signal input
rlabel metal2 s 274822 0 274878 800 6 la_oenb[43]
port 465 nsew signal input
rlabel metal2 s 278134 0 278190 800 6 la_oenb[44]
port 466 nsew signal input
rlabel metal2 s 281446 0 281502 800 6 la_oenb[45]
port 467 nsew signal input
rlabel metal2 s 284758 0 284814 800 6 la_oenb[46]
port 468 nsew signal input
rlabel metal2 s 288070 0 288126 800 6 la_oenb[47]
port 469 nsew signal input
rlabel metal2 s 291382 0 291438 800 6 la_oenb[48]
port 470 nsew signal input
rlabel metal2 s 294694 0 294750 800 6 la_oenb[49]
port 471 nsew signal input
rlabel metal2 s 145654 0 145710 800 6 la_oenb[4]
port 472 nsew signal input
rlabel metal2 s 298006 0 298062 800 6 la_oenb[50]
port 473 nsew signal input
rlabel metal2 s 301318 0 301374 800 6 la_oenb[51]
port 474 nsew signal input
rlabel metal2 s 304630 0 304686 800 6 la_oenb[52]
port 475 nsew signal input
rlabel metal2 s 307942 0 307998 800 6 la_oenb[53]
port 476 nsew signal input
rlabel metal2 s 311254 0 311310 800 6 la_oenb[54]
port 477 nsew signal input
rlabel metal2 s 314566 0 314622 800 6 la_oenb[55]
port 478 nsew signal input
rlabel metal2 s 317878 0 317934 800 6 la_oenb[56]
port 479 nsew signal input
rlabel metal2 s 321190 0 321246 800 6 la_oenb[57]
port 480 nsew signal input
rlabel metal2 s 324502 0 324558 800 6 la_oenb[58]
port 481 nsew signal input
rlabel metal2 s 327814 0 327870 800 6 la_oenb[59]
port 482 nsew signal input
rlabel metal2 s 148966 0 149022 800 6 la_oenb[5]
port 483 nsew signal input
rlabel metal2 s 331126 0 331182 800 6 la_oenb[60]
port 484 nsew signal input
rlabel metal2 s 334438 0 334494 800 6 la_oenb[61]
port 485 nsew signal input
rlabel metal2 s 337750 0 337806 800 6 la_oenb[62]
port 486 nsew signal input
rlabel metal2 s 341062 0 341118 800 6 la_oenb[63]
port 487 nsew signal input
rlabel metal2 s 344374 0 344430 800 6 la_oenb[64]
port 488 nsew signal input
rlabel metal2 s 347686 0 347742 800 6 la_oenb[65]
port 489 nsew signal input
rlabel metal2 s 350998 0 351054 800 6 la_oenb[66]
port 490 nsew signal input
rlabel metal2 s 354310 0 354366 800 6 la_oenb[67]
port 491 nsew signal input
rlabel metal2 s 357622 0 357678 800 6 la_oenb[68]
port 492 nsew signal input
rlabel metal2 s 360934 0 360990 800 6 la_oenb[69]
port 493 nsew signal input
rlabel metal2 s 152278 0 152334 800 6 la_oenb[6]
port 494 nsew signal input
rlabel metal2 s 364246 0 364302 800 6 la_oenb[70]
port 495 nsew signal input
rlabel metal2 s 367558 0 367614 800 6 la_oenb[71]
port 496 nsew signal input
rlabel metal2 s 370870 0 370926 800 6 la_oenb[72]
port 497 nsew signal input
rlabel metal2 s 374182 0 374238 800 6 la_oenb[73]
port 498 nsew signal input
rlabel metal2 s 377494 0 377550 800 6 la_oenb[74]
port 499 nsew signal input
rlabel metal2 s 380806 0 380862 800 6 la_oenb[75]
port 500 nsew signal input
rlabel metal2 s 384118 0 384174 800 6 la_oenb[76]
port 501 nsew signal input
rlabel metal2 s 387430 0 387486 800 6 la_oenb[77]
port 502 nsew signal input
rlabel metal2 s 390742 0 390798 800 6 la_oenb[78]
port 503 nsew signal input
rlabel metal2 s 394054 0 394110 800 6 la_oenb[79]
port 504 nsew signal input
rlabel metal2 s 155590 0 155646 800 6 la_oenb[7]
port 505 nsew signal input
rlabel metal2 s 397366 0 397422 800 6 la_oenb[80]
port 506 nsew signal input
rlabel metal2 s 400678 0 400734 800 6 la_oenb[81]
port 507 nsew signal input
rlabel metal2 s 403990 0 404046 800 6 la_oenb[82]
port 508 nsew signal input
rlabel metal2 s 407302 0 407358 800 6 la_oenb[83]
port 509 nsew signal input
rlabel metal2 s 410614 0 410670 800 6 la_oenb[84]
port 510 nsew signal input
rlabel metal2 s 413926 0 413982 800 6 la_oenb[85]
port 511 nsew signal input
rlabel metal2 s 417238 0 417294 800 6 la_oenb[86]
port 512 nsew signal input
rlabel metal2 s 420550 0 420606 800 6 la_oenb[87]
port 513 nsew signal input
rlabel metal2 s 423862 0 423918 800 6 la_oenb[88]
port 514 nsew signal input
rlabel metal2 s 427174 0 427230 800 6 la_oenb[89]
port 515 nsew signal input
rlabel metal2 s 158902 0 158958 800 6 la_oenb[8]
port 516 nsew signal input
rlabel metal2 s 430486 0 430542 800 6 la_oenb[90]
port 517 nsew signal input
rlabel metal2 s 433798 0 433854 800 6 la_oenb[91]
port 518 nsew signal input
rlabel metal2 s 437110 0 437166 800 6 la_oenb[92]
port 519 nsew signal input
rlabel metal2 s 440422 0 440478 800 6 la_oenb[93]
port 520 nsew signal input
rlabel metal2 s 443734 0 443790 800 6 la_oenb[94]
port 521 nsew signal input
rlabel metal2 s 447046 0 447102 800 6 la_oenb[95]
port 522 nsew signal input
rlabel metal2 s 450358 0 450414 800 6 la_oenb[96]
port 523 nsew signal input
rlabel metal2 s 453670 0 453726 800 6 la_oenb[97]
port 524 nsew signal input
rlabel metal2 s 456982 0 457038 800 6 la_oenb[98]
port 525 nsew signal input
rlabel metal2 s 460294 0 460350 800 6 la_oenb[99]
port 526 nsew signal input
rlabel metal2 s 162214 0 162270 800 6 la_oenb[9]
port 527 nsew signal input
rlabel metal2 s 554134 0 554190 800 6 user_clock2
port 528 nsew signal input
rlabel metal2 s 555238 0 555294 800 6 user_irq[0]
port 529 nsew signal output
rlabel metal2 s 556342 0 556398 800 6 user_irq[1]
port 530 nsew signal output
rlabel metal2 s 557446 0 557502 800 6 user_irq[2]
port 531 nsew signal output
rlabel metal4 s 4208 2128 4528 684400 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 684400 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 684400 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 684400 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 684400 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 684400 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 684400 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 684400 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 684400 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 684400 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 684400 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 684400 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 372848 2128 373168 684400 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 403568 2128 403888 684400 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 434288 2128 434608 684400 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 465008 2128 465328 684400 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 495728 2128 496048 684400 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 526448 2128 526768 684400 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 557168 2128 557488 684400 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 684400 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 684400 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 684400 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 684400 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 684400 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 684400 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 684400 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 684400 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 684400 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 684400 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 684400 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 684400 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 388208 2128 388528 684400 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 418928 2128 419248 684400 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 449648 2128 449968 684400 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 480368 2128 480688 684400 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 511088 2128 511408 684400 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 541808 2128 542128 684400 6 vssd1
port 533 nsew ground bidirectional
rlabel metal2 s 13174 0 13230 800 6 wb_clk_i
port 534 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 wb_rst_i
port 535 nsew signal input
rlabel metal2 s 15382 0 15438 800 6 wbs_ack_o
port 536 nsew signal output
rlabel metal2 s 19798 0 19854 800 6 wbs_adr_i[0]
port 537 nsew signal input
rlabel metal2 s 57334 0 57390 800 6 wbs_adr_i[10]
port 538 nsew signal input
rlabel metal2 s 60646 0 60702 800 6 wbs_adr_i[11]
port 539 nsew signal input
rlabel metal2 s 63958 0 64014 800 6 wbs_adr_i[12]
port 540 nsew signal input
rlabel metal2 s 67270 0 67326 800 6 wbs_adr_i[13]
port 541 nsew signal input
rlabel metal2 s 70582 0 70638 800 6 wbs_adr_i[14]
port 542 nsew signal input
rlabel metal2 s 73894 0 73950 800 6 wbs_adr_i[15]
port 543 nsew signal input
rlabel metal2 s 77206 0 77262 800 6 wbs_adr_i[16]
port 544 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 wbs_adr_i[17]
port 545 nsew signal input
rlabel metal2 s 83830 0 83886 800 6 wbs_adr_i[18]
port 546 nsew signal input
rlabel metal2 s 87142 0 87198 800 6 wbs_adr_i[19]
port 547 nsew signal input
rlabel metal2 s 24214 0 24270 800 6 wbs_adr_i[1]
port 548 nsew signal input
rlabel metal2 s 90454 0 90510 800 6 wbs_adr_i[20]
port 549 nsew signal input
rlabel metal2 s 93766 0 93822 800 6 wbs_adr_i[21]
port 550 nsew signal input
rlabel metal2 s 97078 0 97134 800 6 wbs_adr_i[22]
port 551 nsew signal input
rlabel metal2 s 100390 0 100446 800 6 wbs_adr_i[23]
port 552 nsew signal input
rlabel metal2 s 103702 0 103758 800 6 wbs_adr_i[24]
port 553 nsew signal input
rlabel metal2 s 107014 0 107070 800 6 wbs_adr_i[25]
port 554 nsew signal input
rlabel metal2 s 110326 0 110382 800 6 wbs_adr_i[26]
port 555 nsew signal input
rlabel metal2 s 113638 0 113694 800 6 wbs_adr_i[27]
port 556 nsew signal input
rlabel metal2 s 116950 0 117006 800 6 wbs_adr_i[28]
port 557 nsew signal input
rlabel metal2 s 120262 0 120318 800 6 wbs_adr_i[29]
port 558 nsew signal input
rlabel metal2 s 28630 0 28686 800 6 wbs_adr_i[2]
port 559 nsew signal input
rlabel metal2 s 123574 0 123630 800 6 wbs_adr_i[30]
port 560 nsew signal input
rlabel metal2 s 126886 0 126942 800 6 wbs_adr_i[31]
port 561 nsew signal input
rlabel metal2 s 33046 0 33102 800 6 wbs_adr_i[3]
port 562 nsew signal input
rlabel metal2 s 37462 0 37518 800 6 wbs_adr_i[4]
port 563 nsew signal input
rlabel metal2 s 40774 0 40830 800 6 wbs_adr_i[5]
port 564 nsew signal input
rlabel metal2 s 44086 0 44142 800 6 wbs_adr_i[6]
port 565 nsew signal input
rlabel metal2 s 47398 0 47454 800 6 wbs_adr_i[7]
port 566 nsew signal input
rlabel metal2 s 50710 0 50766 800 6 wbs_adr_i[8]
port 567 nsew signal input
rlabel metal2 s 54022 0 54078 800 6 wbs_adr_i[9]
port 568 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 wbs_cyc_i
port 569 nsew signal input
rlabel metal2 s 20902 0 20958 800 6 wbs_dat_i[0]
port 570 nsew signal input
rlabel metal2 s 58438 0 58494 800 6 wbs_dat_i[10]
port 571 nsew signal input
rlabel metal2 s 61750 0 61806 800 6 wbs_dat_i[11]
port 572 nsew signal input
rlabel metal2 s 65062 0 65118 800 6 wbs_dat_i[12]
port 573 nsew signal input
rlabel metal2 s 68374 0 68430 800 6 wbs_dat_i[13]
port 574 nsew signal input
rlabel metal2 s 71686 0 71742 800 6 wbs_dat_i[14]
port 575 nsew signal input
rlabel metal2 s 74998 0 75054 800 6 wbs_dat_i[15]
port 576 nsew signal input
rlabel metal2 s 78310 0 78366 800 6 wbs_dat_i[16]
port 577 nsew signal input
rlabel metal2 s 81622 0 81678 800 6 wbs_dat_i[17]
port 578 nsew signal input
rlabel metal2 s 84934 0 84990 800 6 wbs_dat_i[18]
port 579 nsew signal input
rlabel metal2 s 88246 0 88302 800 6 wbs_dat_i[19]
port 580 nsew signal input
rlabel metal2 s 25318 0 25374 800 6 wbs_dat_i[1]
port 581 nsew signal input
rlabel metal2 s 91558 0 91614 800 6 wbs_dat_i[20]
port 582 nsew signal input
rlabel metal2 s 94870 0 94926 800 6 wbs_dat_i[21]
port 583 nsew signal input
rlabel metal2 s 98182 0 98238 800 6 wbs_dat_i[22]
port 584 nsew signal input
rlabel metal2 s 101494 0 101550 800 6 wbs_dat_i[23]
port 585 nsew signal input
rlabel metal2 s 104806 0 104862 800 6 wbs_dat_i[24]
port 586 nsew signal input
rlabel metal2 s 108118 0 108174 800 6 wbs_dat_i[25]
port 587 nsew signal input
rlabel metal2 s 111430 0 111486 800 6 wbs_dat_i[26]
port 588 nsew signal input
rlabel metal2 s 114742 0 114798 800 6 wbs_dat_i[27]
port 589 nsew signal input
rlabel metal2 s 118054 0 118110 800 6 wbs_dat_i[28]
port 590 nsew signal input
rlabel metal2 s 121366 0 121422 800 6 wbs_dat_i[29]
port 591 nsew signal input
rlabel metal2 s 29734 0 29790 800 6 wbs_dat_i[2]
port 592 nsew signal input
rlabel metal2 s 124678 0 124734 800 6 wbs_dat_i[30]
port 593 nsew signal input
rlabel metal2 s 127990 0 128046 800 6 wbs_dat_i[31]
port 594 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 wbs_dat_i[3]
port 595 nsew signal input
rlabel metal2 s 38566 0 38622 800 6 wbs_dat_i[4]
port 596 nsew signal input
rlabel metal2 s 41878 0 41934 800 6 wbs_dat_i[5]
port 597 nsew signal input
rlabel metal2 s 45190 0 45246 800 6 wbs_dat_i[6]
port 598 nsew signal input
rlabel metal2 s 48502 0 48558 800 6 wbs_dat_i[7]
port 599 nsew signal input
rlabel metal2 s 51814 0 51870 800 6 wbs_dat_i[8]
port 600 nsew signal input
rlabel metal2 s 55126 0 55182 800 6 wbs_dat_i[9]
port 601 nsew signal input
rlabel metal2 s 22006 0 22062 800 6 wbs_dat_o[0]
port 602 nsew signal output
rlabel metal2 s 59542 0 59598 800 6 wbs_dat_o[10]
port 603 nsew signal output
rlabel metal2 s 62854 0 62910 800 6 wbs_dat_o[11]
port 604 nsew signal output
rlabel metal2 s 66166 0 66222 800 6 wbs_dat_o[12]
port 605 nsew signal output
rlabel metal2 s 69478 0 69534 800 6 wbs_dat_o[13]
port 606 nsew signal output
rlabel metal2 s 72790 0 72846 800 6 wbs_dat_o[14]
port 607 nsew signal output
rlabel metal2 s 76102 0 76158 800 6 wbs_dat_o[15]
port 608 nsew signal output
rlabel metal2 s 79414 0 79470 800 6 wbs_dat_o[16]
port 609 nsew signal output
rlabel metal2 s 82726 0 82782 800 6 wbs_dat_o[17]
port 610 nsew signal output
rlabel metal2 s 86038 0 86094 800 6 wbs_dat_o[18]
port 611 nsew signal output
rlabel metal2 s 89350 0 89406 800 6 wbs_dat_o[19]
port 612 nsew signal output
rlabel metal2 s 26422 0 26478 800 6 wbs_dat_o[1]
port 613 nsew signal output
rlabel metal2 s 92662 0 92718 800 6 wbs_dat_o[20]
port 614 nsew signal output
rlabel metal2 s 95974 0 96030 800 6 wbs_dat_o[21]
port 615 nsew signal output
rlabel metal2 s 99286 0 99342 800 6 wbs_dat_o[22]
port 616 nsew signal output
rlabel metal2 s 102598 0 102654 800 6 wbs_dat_o[23]
port 617 nsew signal output
rlabel metal2 s 105910 0 105966 800 6 wbs_dat_o[24]
port 618 nsew signal output
rlabel metal2 s 109222 0 109278 800 6 wbs_dat_o[25]
port 619 nsew signal output
rlabel metal2 s 112534 0 112590 800 6 wbs_dat_o[26]
port 620 nsew signal output
rlabel metal2 s 115846 0 115902 800 6 wbs_dat_o[27]
port 621 nsew signal output
rlabel metal2 s 119158 0 119214 800 6 wbs_dat_o[28]
port 622 nsew signal output
rlabel metal2 s 122470 0 122526 800 6 wbs_dat_o[29]
port 623 nsew signal output
rlabel metal2 s 30838 0 30894 800 6 wbs_dat_o[2]
port 624 nsew signal output
rlabel metal2 s 125782 0 125838 800 6 wbs_dat_o[30]
port 625 nsew signal output
rlabel metal2 s 129094 0 129150 800 6 wbs_dat_o[31]
port 626 nsew signal output
rlabel metal2 s 35254 0 35310 800 6 wbs_dat_o[3]
port 627 nsew signal output
rlabel metal2 s 39670 0 39726 800 6 wbs_dat_o[4]
port 628 nsew signal output
rlabel metal2 s 42982 0 43038 800 6 wbs_dat_o[5]
port 629 nsew signal output
rlabel metal2 s 46294 0 46350 800 6 wbs_dat_o[6]
port 630 nsew signal output
rlabel metal2 s 49606 0 49662 800 6 wbs_dat_o[7]
port 631 nsew signal output
rlabel metal2 s 52918 0 52974 800 6 wbs_dat_o[8]
port 632 nsew signal output
rlabel metal2 s 56230 0 56286 800 6 wbs_dat_o[9]
port 633 nsew signal output
rlabel metal2 s 23110 0 23166 800 6 wbs_sel_i[0]
port 634 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 wbs_sel_i[1]
port 635 nsew signal input
rlabel metal2 s 31942 0 31998 800 6 wbs_sel_i[2]
port 636 nsew signal input
rlabel metal2 s 36358 0 36414 800 6 wbs_sel_i[3]
port 637 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 wbs_stb_i
port 638 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 wbs_we_i
port 639 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 570805 686669
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 995002590
string GDS_FILE /mnt/r/work/Rift2Go_2330_Sky130_MPW8/openlane/user_proj_example/runs/22_12_29_15_16/results/signoff/rift2Wrap.magic.gds
string GDS_START 2025804
<< end >>

