VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO rift2Wrap
  CLASS BLOCK ;
  FOREIGN rift2Wrap ;
  ORIGIN 0.000 0.000 ;
  SIZE 2854.025 BY 3433.345 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 1393.360 2854.025 1393.960 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2178.190 3429.345 2178.470 3433.345 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1861.710 3429.345 1861.990 3433.345 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1545.230 3429.345 1545.510 3433.345 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1228.750 3429.345 1229.030 3433.345 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 912.270 3429.345 912.550 3433.345 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.790 3429.345 596.070 3433.345 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.310 3429.345 279.590 3433.345 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3391.880 4.000 3392.480 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3138.920 4.000 3139.520 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2885.960 4.000 2886.560 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 1651.760 2854.025 1652.360 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2633.000 4.000 2633.600 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2380.040 4.000 2380.640 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2127.080 4.000 2127.680 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1874.120 4.000 1874.720 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1621.160 4.000 1621.760 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1368.200 4.000 1368.800 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1115.240 4.000 1115.840 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 862.280 4.000 862.880 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 609.320 4.000 609.920 ;
    END
  END analog_io[28]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 1910.160 2854.025 1910.760 ;
    END
  END analog_io[2]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 2168.560 2854.025 2169.160 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 2426.960 2854.025 2427.560 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 2685.360 2854.025 2685.960 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 2943.760 2854.025 2944.360 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 3202.160 2854.025 3202.760 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2811.150 3429.345 2811.430 3433.345 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2494.670 3429.345 2494.950 3433.345 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 36.760 2854.025 37.360 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 2233.160 2854.025 2233.760 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 2491.560 2854.025 2492.160 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 2749.960 2854.025 2750.560 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 3008.360 2854.025 3008.960 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 3266.760 2854.025 3267.360 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2732.030 3429.345 2732.310 3433.345 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2415.550 3429.345 2415.830 3433.345 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2099.070 3429.345 2099.350 3433.345 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1782.590 3429.345 1782.870 3433.345 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1466.110 3429.345 1466.390 3433.345 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 230.560 2854.025 231.160 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1149.630 3429.345 1149.910 3433.345 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 833.150 3429.345 833.430 3433.345 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.670 3429.345 516.950 3433.345 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 3429.345 200.470 3433.345 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3328.640 4.000 3329.240 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3075.680 4.000 3076.280 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2822.720 4.000 2823.320 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2569.760 4.000 2570.360 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2316.800 4.000 2317.400 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2063.840 4.000 2064.440 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 424.360 2854.025 424.960 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1810.880 4.000 1811.480 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1557.920 4.000 1558.520 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1304.960 4.000 1305.560 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1052.000 4.000 1052.600 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 799.040 4.000 799.640 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 546.080 4.000 546.680 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 356.360 4.000 356.960 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 618.160 2854.025 618.760 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 811.960 2854.025 812.560 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 1005.760 2854.025 1006.360 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 1199.560 2854.025 1200.160 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 1457.960 2854.025 1458.560 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 1716.360 2854.025 1716.960 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 1974.760 2854.025 1975.360 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 165.960 2854.025 166.560 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 2362.360 2854.025 2362.960 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 2620.760 2854.025 2621.360 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 2879.160 2854.025 2879.760 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 3137.560 2854.025 3138.160 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 3395.960 2854.025 3396.560 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2573.790 3429.345 2574.070 3433.345 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2257.310 3429.345 2257.590 3433.345 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1940.830 3429.345 1941.110 3433.345 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1624.350 3429.345 1624.630 3433.345 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1307.870 3429.345 1308.150 3433.345 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 359.760 2854.025 360.360 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 991.390 3429.345 991.670 3433.345 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.910 3429.345 675.190 3433.345 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.430 3429.345 358.710 3433.345 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 3429.345 42.230 3433.345 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3202.160 4.000 3202.760 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2949.200 4.000 2949.800 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2696.240 4.000 2696.840 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2443.280 4.000 2443.880 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2190.320 4.000 2190.920 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1937.360 4.000 1937.960 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 553.560 2854.025 554.160 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1684.400 4.000 1685.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1431.440 4.000 1432.040 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1178.480 4.000 1179.080 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 925.520 4.000 926.120 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 672.560 4.000 673.160 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 419.600 4.000 420.200 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.880 4.000 230.480 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.160 4.000 40.760 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 747.360 2854.025 747.960 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 941.160 2854.025 941.760 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 1134.960 2854.025 1135.560 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 1328.760 2854.025 1329.360 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 1587.160 2854.025 1587.760 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 1845.560 2854.025 1846.160 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 2103.960 2854.025 2104.560 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 101.360 2854.025 101.960 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 2297.760 2854.025 2298.360 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 2556.160 2854.025 2556.760 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 2814.560 2854.025 2815.160 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 3072.960 2854.025 3073.560 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 3331.360 2854.025 3331.960 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2652.910 3429.345 2653.190 3433.345 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2336.430 3429.345 2336.710 3433.345 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2019.950 3429.345 2020.230 3433.345 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1703.470 3429.345 1703.750 3433.345 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1386.990 3429.345 1387.270 3433.345 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 295.160 2854.025 295.760 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1070.510 3429.345 1070.790 3433.345 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.030 3429.345 754.310 3433.345 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.550 3429.345 437.830 3433.345 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.070 3429.345 121.350 3433.345 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3265.400 4.000 3266.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3012.440 4.000 3013.040 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2759.480 4.000 2760.080 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2506.520 4.000 2507.120 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2253.560 4.000 2254.160 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2000.600 4.000 2001.200 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 488.960 2854.025 489.560 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1747.640 4.000 1748.240 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1494.680 4.000 1495.280 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1241.720 4.000 1242.320 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 988.760 4.000 989.360 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 735.800 4.000 736.400 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.840 4.000 483.440 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.120 4.000 293.720 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 4.000 104.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 682.760 2854.025 683.360 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 876.560 2854.025 877.160 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 1070.360 2854.025 1070.960 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 1264.160 2854.025 1264.760 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 1522.560 2854.025 1523.160 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 1780.960 2854.025 1781.560 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2850.025 2039.360 2854.025 2039.960 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.990 0.000 651.270 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2306.990 0.000 2307.270 4.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2323.550 0.000 2323.830 4.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2340.110 0.000 2340.390 4.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2356.670 0.000 2356.950 4.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2373.230 0.000 2373.510 4.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2389.790 0.000 2390.070 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2406.350 0.000 2406.630 4.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2422.910 0.000 2423.190 4.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2439.470 0.000 2439.750 4.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2456.030 0.000 2456.310 4.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 816.590 0.000 816.870 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2472.590 0.000 2472.870 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2489.150 0.000 2489.430 4.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2505.710 0.000 2505.990 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2522.270 0.000 2522.550 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2538.830 0.000 2539.110 4.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2555.390 0.000 2555.670 4.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2571.950 0.000 2572.230 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2588.510 0.000 2588.790 4.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2605.070 0.000 2605.350 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2621.630 0.000 2621.910 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 833.150 0.000 833.430 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2638.190 0.000 2638.470 4.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2654.750 0.000 2655.030 4.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2671.310 0.000 2671.590 4.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2687.870 0.000 2688.150 4.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2704.430 0.000 2704.710 4.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2720.990 0.000 2721.270 4.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2737.550 0.000 2737.830 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2754.110 0.000 2754.390 4.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 849.710 0.000 849.990 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 866.270 0.000 866.550 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.830 0.000 883.110 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 899.390 0.000 899.670 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.950 0.000 916.230 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.510 0.000 932.790 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.070 0.000 949.350 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 965.630 0.000 965.910 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.550 0.000 667.830 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 982.190 0.000 982.470 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.750 0.000 999.030 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1015.310 0.000 1015.590 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1031.870 0.000 1032.150 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1048.430 0.000 1048.710 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1064.990 0.000 1065.270 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1081.550 0.000 1081.830 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1098.110 0.000 1098.390 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1114.670 0.000 1114.950 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1131.230 0.000 1131.510 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 684.110 0.000 684.390 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1147.790 0.000 1148.070 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1164.350 0.000 1164.630 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1180.910 0.000 1181.190 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1197.470 0.000 1197.750 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1214.030 0.000 1214.310 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1230.590 0.000 1230.870 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1247.150 0.000 1247.430 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1263.710 0.000 1263.990 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1280.270 0.000 1280.550 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1296.830 0.000 1297.110 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.670 0.000 700.950 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1313.390 0.000 1313.670 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1329.950 0.000 1330.230 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1346.510 0.000 1346.790 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1363.070 0.000 1363.350 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1379.630 0.000 1379.910 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1396.190 0.000 1396.470 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1412.750 0.000 1413.030 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1429.310 0.000 1429.590 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1445.870 0.000 1446.150 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1462.430 0.000 1462.710 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.230 0.000 717.510 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1478.990 0.000 1479.270 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1495.550 0.000 1495.830 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1512.110 0.000 1512.390 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1528.670 0.000 1528.950 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1545.230 0.000 1545.510 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1561.790 0.000 1562.070 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1578.350 0.000 1578.630 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1594.910 0.000 1595.190 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1611.470 0.000 1611.750 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1628.030 0.000 1628.310 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 733.790 0.000 734.070 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1644.590 0.000 1644.870 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1661.150 0.000 1661.430 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1677.710 0.000 1677.990 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1694.270 0.000 1694.550 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1710.830 0.000 1711.110 4.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1727.390 0.000 1727.670 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1743.950 0.000 1744.230 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1760.510 0.000 1760.790 4.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1777.070 0.000 1777.350 4.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1793.630 0.000 1793.910 4.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.350 0.000 750.630 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1810.190 0.000 1810.470 4.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1826.750 0.000 1827.030 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1843.310 0.000 1843.590 4.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1859.870 0.000 1860.150 4.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1876.430 0.000 1876.710 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1892.990 0.000 1893.270 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1909.550 0.000 1909.830 4.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1926.110 0.000 1926.390 4.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1942.670 0.000 1942.950 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1959.230 0.000 1959.510 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.910 0.000 767.190 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1975.790 0.000 1976.070 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1992.350 0.000 1992.630 4.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2008.910 0.000 2009.190 4.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2025.470 0.000 2025.750 4.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2042.030 0.000 2042.310 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2058.590 0.000 2058.870 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2075.150 0.000 2075.430 4.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2091.710 0.000 2091.990 4.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2108.270 0.000 2108.550 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2124.830 0.000 2125.110 4.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.470 0.000 783.750 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2141.390 0.000 2141.670 4.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2157.950 0.000 2158.230 4.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2174.510 0.000 2174.790 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2191.070 0.000 2191.350 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2207.630 0.000 2207.910 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2224.190 0.000 2224.470 4.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2240.750 0.000 2241.030 4.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2257.310 0.000 2257.590 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2273.870 0.000 2274.150 4.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2290.430 0.000 2290.710 4.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.030 0.000 800.310 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.510 0.000 656.790 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2312.510 0.000 2312.790 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2329.070 0.000 2329.350 4.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2345.630 0.000 2345.910 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2362.190 0.000 2362.470 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2378.750 0.000 2379.030 4.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2395.310 0.000 2395.590 4.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2411.870 0.000 2412.150 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2428.430 0.000 2428.710 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2444.990 0.000 2445.270 4.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2461.550 0.000 2461.830 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 822.110 0.000 822.390 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2478.110 0.000 2478.390 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2494.670 0.000 2494.950 4.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2511.230 0.000 2511.510 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2527.790 0.000 2528.070 4.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2544.350 0.000 2544.630 4.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2560.910 0.000 2561.190 4.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2577.470 0.000 2577.750 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2594.030 0.000 2594.310 4.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2610.590 0.000 2610.870 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2627.150 0.000 2627.430 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 838.670 0.000 838.950 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2643.710 0.000 2643.990 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2660.270 0.000 2660.550 4.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2676.830 0.000 2677.110 4.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2693.390 0.000 2693.670 4.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2709.950 0.000 2710.230 4.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2726.510 0.000 2726.790 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2743.070 0.000 2743.350 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2759.630 0.000 2759.910 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 855.230 0.000 855.510 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.790 0.000 872.070 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.350 0.000 888.630 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 904.910 0.000 905.190 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.470 0.000 921.750 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 938.030 0.000 938.310 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 954.590 0.000 954.870 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 971.150 0.000 971.430 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.070 0.000 673.350 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 987.710 0.000 987.990 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1004.270 0.000 1004.550 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1020.830 0.000 1021.110 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1037.390 0.000 1037.670 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1053.950 0.000 1054.230 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1070.510 0.000 1070.790 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1087.070 0.000 1087.350 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1103.630 0.000 1103.910 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1120.190 0.000 1120.470 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1136.750 0.000 1137.030 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.630 0.000 689.910 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1153.310 0.000 1153.590 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1169.870 0.000 1170.150 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1186.430 0.000 1186.710 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1202.990 0.000 1203.270 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1219.550 0.000 1219.830 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1236.110 0.000 1236.390 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1252.670 0.000 1252.950 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1269.230 0.000 1269.510 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1285.790 0.000 1286.070 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1302.350 0.000 1302.630 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.190 0.000 706.470 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1318.910 0.000 1319.190 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1335.470 0.000 1335.750 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1352.030 0.000 1352.310 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1368.590 0.000 1368.870 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1385.150 0.000 1385.430 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1401.710 0.000 1401.990 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1418.270 0.000 1418.550 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1434.830 0.000 1435.110 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1451.390 0.000 1451.670 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1467.950 0.000 1468.230 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.750 0.000 723.030 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1484.510 0.000 1484.790 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1501.070 0.000 1501.350 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1517.630 0.000 1517.910 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1534.190 0.000 1534.470 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1550.750 0.000 1551.030 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1567.310 0.000 1567.590 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1583.870 0.000 1584.150 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1600.430 0.000 1600.710 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1616.990 0.000 1617.270 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1633.550 0.000 1633.830 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 739.310 0.000 739.590 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1650.110 0.000 1650.390 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1666.670 0.000 1666.950 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1683.230 0.000 1683.510 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1699.790 0.000 1700.070 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1716.350 0.000 1716.630 4.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1732.910 0.000 1733.190 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1749.470 0.000 1749.750 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1766.030 0.000 1766.310 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1782.590 0.000 1782.870 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1799.150 0.000 1799.430 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 755.870 0.000 756.150 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1815.710 0.000 1815.990 4.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1832.270 0.000 1832.550 4.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1848.830 0.000 1849.110 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1865.390 0.000 1865.670 4.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1881.950 0.000 1882.230 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1898.510 0.000 1898.790 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1915.070 0.000 1915.350 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1931.630 0.000 1931.910 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1948.190 0.000 1948.470 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1964.750 0.000 1965.030 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.430 0.000 772.710 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1981.310 0.000 1981.590 4.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1997.870 0.000 1998.150 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2014.430 0.000 2014.710 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2030.990 0.000 2031.270 4.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2047.550 0.000 2047.830 4.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2064.110 0.000 2064.390 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2080.670 0.000 2080.950 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2097.230 0.000 2097.510 4.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2113.790 0.000 2114.070 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2130.350 0.000 2130.630 4.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.990 0.000 789.270 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2146.910 0.000 2147.190 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2163.470 0.000 2163.750 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2180.030 0.000 2180.310 4.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2196.590 0.000 2196.870 4.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2213.150 0.000 2213.430 4.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2229.710 0.000 2229.990 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2246.270 0.000 2246.550 4.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2262.830 0.000 2263.110 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2279.390 0.000 2279.670 4.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2295.950 0.000 2296.230 4.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.550 0.000 805.830 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.030 0.000 662.310 4.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2318.030 0.000 2318.310 4.000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2334.590 0.000 2334.870 4.000 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2351.150 0.000 2351.430 4.000 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2367.710 0.000 2367.990 4.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2384.270 0.000 2384.550 4.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2400.830 0.000 2401.110 4.000 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2417.390 0.000 2417.670 4.000 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2433.950 0.000 2434.230 4.000 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2450.510 0.000 2450.790 4.000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2467.070 0.000 2467.350 4.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 827.630 0.000 827.910 4.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2483.630 0.000 2483.910 4.000 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2500.190 0.000 2500.470 4.000 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2516.750 0.000 2517.030 4.000 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2533.310 0.000 2533.590 4.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2549.870 0.000 2550.150 4.000 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2566.430 0.000 2566.710 4.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2582.990 0.000 2583.270 4.000 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2599.550 0.000 2599.830 4.000 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2616.110 0.000 2616.390 4.000 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2632.670 0.000 2632.950 4.000 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 844.190 0.000 844.470 4.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2649.230 0.000 2649.510 4.000 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2665.790 0.000 2666.070 4.000 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2682.350 0.000 2682.630 4.000 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2698.910 0.000 2699.190 4.000 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2715.470 0.000 2715.750 4.000 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2732.030 0.000 2732.310 4.000 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2748.590 0.000 2748.870 4.000 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2765.150 0.000 2765.430 4.000 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 860.750 0.000 861.030 4.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.310 0.000 877.590 4.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 893.870 0.000 894.150 4.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 910.430 0.000 910.710 4.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 926.990 0.000 927.270 4.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 943.550 0.000 943.830 4.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 960.110 0.000 960.390 4.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 976.670 0.000 976.950 4.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 678.590 0.000 678.870 4.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 993.230 0.000 993.510 4.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1009.790 0.000 1010.070 4.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1026.350 0.000 1026.630 4.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1042.910 0.000 1043.190 4.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.470 0.000 1059.750 4.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1076.030 0.000 1076.310 4.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1092.590 0.000 1092.870 4.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1109.150 0.000 1109.430 4.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1125.710 0.000 1125.990 4.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1142.270 0.000 1142.550 4.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.150 0.000 695.430 4.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1158.830 0.000 1159.110 4.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.390 0.000 1175.670 4.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1191.950 0.000 1192.230 4.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1208.510 0.000 1208.790 4.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1225.070 0.000 1225.350 4.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1241.630 0.000 1241.910 4.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1258.190 0.000 1258.470 4.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1274.750 0.000 1275.030 4.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.310 0.000 1291.590 4.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1307.870 0.000 1308.150 4.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.710 0.000 711.990 4.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1324.430 0.000 1324.710 4.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1340.990 0.000 1341.270 4.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1357.550 0.000 1357.830 4.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1374.110 0.000 1374.390 4.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1390.670 0.000 1390.950 4.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1407.230 0.000 1407.510 4.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1423.790 0.000 1424.070 4.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1440.350 0.000 1440.630 4.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1456.910 0.000 1457.190 4.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1473.470 0.000 1473.750 4.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.270 0.000 728.550 4.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1490.030 0.000 1490.310 4.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1506.590 0.000 1506.870 4.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1523.150 0.000 1523.430 4.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1539.710 0.000 1539.990 4.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1556.270 0.000 1556.550 4.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1572.830 0.000 1573.110 4.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1589.390 0.000 1589.670 4.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1605.950 0.000 1606.230 4.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1622.510 0.000 1622.790 4.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1639.070 0.000 1639.350 4.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 744.830 0.000 745.110 4.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1655.630 0.000 1655.910 4.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1672.190 0.000 1672.470 4.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1688.750 0.000 1689.030 4.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1705.310 0.000 1705.590 4.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1721.870 0.000 1722.150 4.000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1738.430 0.000 1738.710 4.000 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1754.990 0.000 1755.270 4.000 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1771.550 0.000 1771.830 4.000 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1788.110 0.000 1788.390 4.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1804.670 0.000 1804.950 4.000 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.390 0.000 761.670 4.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1821.230 0.000 1821.510 4.000 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1837.790 0.000 1838.070 4.000 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1854.350 0.000 1854.630 4.000 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1870.910 0.000 1871.190 4.000 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1887.470 0.000 1887.750 4.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1904.030 0.000 1904.310 4.000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1920.590 0.000 1920.870 4.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1937.150 0.000 1937.430 4.000 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1953.710 0.000 1953.990 4.000 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1970.270 0.000 1970.550 4.000 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.950 0.000 778.230 4.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1986.830 0.000 1987.110 4.000 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2003.390 0.000 2003.670 4.000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2019.950 0.000 2020.230 4.000 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2036.510 0.000 2036.790 4.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2053.070 0.000 2053.350 4.000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2069.630 0.000 2069.910 4.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2086.190 0.000 2086.470 4.000 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2102.750 0.000 2103.030 4.000 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2119.310 0.000 2119.590 4.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2135.870 0.000 2136.150 4.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.510 0.000 794.790 4.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2152.430 0.000 2152.710 4.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2168.990 0.000 2169.270 4.000 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2185.550 0.000 2185.830 4.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2202.110 0.000 2202.390 4.000 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2218.670 0.000 2218.950 4.000 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2235.230 0.000 2235.510 4.000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2251.790 0.000 2252.070 4.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2268.350 0.000 2268.630 4.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2284.910 0.000 2285.190 4.000 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2301.470 0.000 2301.750 4.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.070 0.000 811.350 4.000 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2770.670 0.000 2770.950 4.000 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2776.190 0.000 2776.470 4.000 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2781.710 0.000 2781.990 4.000 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2787.230 0.000 2787.510 4.000 ;
    END
  END user_irq[2]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 3422.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 3422.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 3422.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 3422.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 3422.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 3422.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 3422.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 3422.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 3422.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 3422.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 3422.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 3422.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.240 10.640 1865.840 3422.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.840 10.640 2019.440 3422.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2171.440 10.640 2173.040 3422.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2325.040 10.640 2326.640 3422.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2478.640 10.640 2480.240 3422.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2632.240 10.640 2633.840 3422.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2785.840 10.640 2787.440 3422.000 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 3422.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 3422.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 3422.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 3422.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 3422.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 3422.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 3422.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 3422.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 3422.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 3422.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 3422.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1787.440 10.640 1789.040 3422.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1941.040 10.640 1942.640 3422.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2094.640 10.640 2096.240 3422.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2248.240 10.640 2249.840 3422.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2401.840 10.640 2403.440 3422.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2555.440 10.640 2557.040 3422.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2709.040 10.640 2710.640 3422.000 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 0.000 66.150 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 0.000 71.670 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.910 0.000 77.190 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.990 0.000 99.270 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.230 0.000 303.510 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.790 0.000 320.070 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.350 0.000 336.630 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.910 0.000 353.190 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.470 0.000 369.750 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.030 0.000 386.310 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 0.000 402.870 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.150 0.000 419.430 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.710 0.000 435.990 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.070 0.000 121.350 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.270 0.000 452.550 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.830 0.000 469.110 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.390 0.000 485.670 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.950 0.000 502.230 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.510 0.000 518.790 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.070 0.000 535.350 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.630 0.000 551.910 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 568.190 0.000 568.470 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.750 0.000 585.030 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 601.310 0.000 601.590 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.150 0.000 143.430 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.870 0.000 618.150 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.430 0.000 634.710 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.230 0.000 165.510 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.310 0.000 187.590 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.870 0.000 204.150 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.430 0.000 220.710 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.990 0.000 237.270 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.550 0.000 253.830 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.110 0.000 270.390 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 0.000 82.710 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.510 0.000 104.790 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.190 0.000 292.470 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.750 0.000 309.030 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 0.000 325.590 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.870 0.000 342.150 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.430 0.000 358.710 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.990 0.000 375.270 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.550 0.000 391.830 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.110 0.000 408.390 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.670 0.000 424.950 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230 0.000 441.510 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 0.000 126.870 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.790 0.000 458.070 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.350 0.000 474.630 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.910 0.000 491.190 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.470 0.000 507.750 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.030 0.000 524.310 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.590 0.000 540.870 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.150 0.000 557.430 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.710 0.000 573.990 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 590.270 0.000 590.550 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.830 0.000 607.110 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.670 0.000 148.950 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.390 0.000 623.670 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.950 0.000 640.230 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.830 0.000 193.110 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.950 0.000 226.230 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.510 0.000 242.790 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.070 0.000 259.350 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.630 0.000 275.910 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.030 0.000 110.310 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.710 0.000 297.990 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.270 0.000 314.550 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.830 0.000 331.110 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.390 0.000 347.670 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 0.000 364.230 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.510 0.000 380.790 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.070 0.000 397.350 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.630 0.000 413.910 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.190 0.000 430.470 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.750 0.000 447.030 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.310 0.000 463.590 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.870 0.000 480.150 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.430 0.000 496.710 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.990 0.000 513.270 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.550 0.000 529.830 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.110 0.000 546.390 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.670 0.000 562.950 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.230 0.000 579.510 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.790 0.000 596.070 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.350 0.000 612.630 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.190 0.000 154.470 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.910 0.000 629.190 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.470 0.000 645.750 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.270 0.000 176.550 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.350 0.000 198.630 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.910 0.000 215.190 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.470 0.000 231.750 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 0.000 248.310 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.590 0.000 264.870 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.150 0.000 281.430 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.550 0.000 115.830 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.630 0.000 137.910 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.710 0.000 159.990 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.790 0.000 182.070 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 0.000 88.230 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2848.320 3421.845 ;
      LAYER met1 ;
        RECT 1.910 10.640 2853.770 3422.000 ;
      LAYER met2 ;
        RECT 1.930 3429.065 41.670 3429.345 ;
        RECT 42.510 3429.065 120.790 3429.345 ;
        RECT 121.630 3429.065 199.910 3429.345 ;
        RECT 200.750 3429.065 279.030 3429.345 ;
        RECT 279.870 3429.065 358.150 3429.345 ;
        RECT 358.990 3429.065 437.270 3429.345 ;
        RECT 438.110 3429.065 516.390 3429.345 ;
        RECT 517.230 3429.065 595.510 3429.345 ;
        RECT 596.350 3429.065 674.630 3429.345 ;
        RECT 675.470 3429.065 753.750 3429.345 ;
        RECT 754.590 3429.065 832.870 3429.345 ;
        RECT 833.710 3429.065 911.990 3429.345 ;
        RECT 912.830 3429.065 991.110 3429.345 ;
        RECT 991.950 3429.065 1070.230 3429.345 ;
        RECT 1071.070 3429.065 1149.350 3429.345 ;
        RECT 1150.190 3429.065 1228.470 3429.345 ;
        RECT 1229.310 3429.065 1307.590 3429.345 ;
        RECT 1308.430 3429.065 1386.710 3429.345 ;
        RECT 1387.550 3429.065 1465.830 3429.345 ;
        RECT 1466.670 3429.065 1544.950 3429.345 ;
        RECT 1545.790 3429.065 1624.070 3429.345 ;
        RECT 1624.910 3429.065 1703.190 3429.345 ;
        RECT 1704.030 3429.065 1782.310 3429.345 ;
        RECT 1783.150 3429.065 1861.430 3429.345 ;
        RECT 1862.270 3429.065 1940.550 3429.345 ;
        RECT 1941.390 3429.065 2019.670 3429.345 ;
        RECT 2020.510 3429.065 2098.790 3429.345 ;
        RECT 2099.630 3429.065 2177.910 3429.345 ;
        RECT 2178.750 3429.065 2257.030 3429.345 ;
        RECT 2257.870 3429.065 2336.150 3429.345 ;
        RECT 2336.990 3429.065 2415.270 3429.345 ;
        RECT 2416.110 3429.065 2494.390 3429.345 ;
        RECT 2495.230 3429.065 2573.510 3429.345 ;
        RECT 2574.350 3429.065 2652.630 3429.345 ;
        RECT 2653.470 3429.065 2731.750 3429.345 ;
        RECT 2732.590 3429.065 2810.870 3429.345 ;
        RECT 2811.710 3429.065 2853.740 3429.345 ;
        RECT 1.930 4.280 2853.740 3429.065 ;
        RECT 1.930 3.670 65.590 4.280 ;
        RECT 66.430 3.670 71.110 4.280 ;
        RECT 71.950 3.670 76.630 4.280 ;
        RECT 77.470 3.670 82.150 4.280 ;
        RECT 82.990 3.670 87.670 4.280 ;
        RECT 88.510 3.670 93.190 4.280 ;
        RECT 94.030 3.670 98.710 4.280 ;
        RECT 99.550 3.670 104.230 4.280 ;
        RECT 105.070 3.670 109.750 4.280 ;
        RECT 110.590 3.670 115.270 4.280 ;
        RECT 116.110 3.670 120.790 4.280 ;
        RECT 121.630 3.670 126.310 4.280 ;
        RECT 127.150 3.670 131.830 4.280 ;
        RECT 132.670 3.670 137.350 4.280 ;
        RECT 138.190 3.670 142.870 4.280 ;
        RECT 143.710 3.670 148.390 4.280 ;
        RECT 149.230 3.670 153.910 4.280 ;
        RECT 154.750 3.670 159.430 4.280 ;
        RECT 160.270 3.670 164.950 4.280 ;
        RECT 165.790 3.670 170.470 4.280 ;
        RECT 171.310 3.670 175.990 4.280 ;
        RECT 176.830 3.670 181.510 4.280 ;
        RECT 182.350 3.670 187.030 4.280 ;
        RECT 187.870 3.670 192.550 4.280 ;
        RECT 193.390 3.670 198.070 4.280 ;
        RECT 198.910 3.670 203.590 4.280 ;
        RECT 204.430 3.670 209.110 4.280 ;
        RECT 209.950 3.670 214.630 4.280 ;
        RECT 215.470 3.670 220.150 4.280 ;
        RECT 220.990 3.670 225.670 4.280 ;
        RECT 226.510 3.670 231.190 4.280 ;
        RECT 232.030 3.670 236.710 4.280 ;
        RECT 237.550 3.670 242.230 4.280 ;
        RECT 243.070 3.670 247.750 4.280 ;
        RECT 248.590 3.670 253.270 4.280 ;
        RECT 254.110 3.670 258.790 4.280 ;
        RECT 259.630 3.670 264.310 4.280 ;
        RECT 265.150 3.670 269.830 4.280 ;
        RECT 270.670 3.670 275.350 4.280 ;
        RECT 276.190 3.670 280.870 4.280 ;
        RECT 281.710 3.670 286.390 4.280 ;
        RECT 287.230 3.670 291.910 4.280 ;
        RECT 292.750 3.670 297.430 4.280 ;
        RECT 298.270 3.670 302.950 4.280 ;
        RECT 303.790 3.670 308.470 4.280 ;
        RECT 309.310 3.670 313.990 4.280 ;
        RECT 314.830 3.670 319.510 4.280 ;
        RECT 320.350 3.670 325.030 4.280 ;
        RECT 325.870 3.670 330.550 4.280 ;
        RECT 331.390 3.670 336.070 4.280 ;
        RECT 336.910 3.670 341.590 4.280 ;
        RECT 342.430 3.670 347.110 4.280 ;
        RECT 347.950 3.670 352.630 4.280 ;
        RECT 353.470 3.670 358.150 4.280 ;
        RECT 358.990 3.670 363.670 4.280 ;
        RECT 364.510 3.670 369.190 4.280 ;
        RECT 370.030 3.670 374.710 4.280 ;
        RECT 375.550 3.670 380.230 4.280 ;
        RECT 381.070 3.670 385.750 4.280 ;
        RECT 386.590 3.670 391.270 4.280 ;
        RECT 392.110 3.670 396.790 4.280 ;
        RECT 397.630 3.670 402.310 4.280 ;
        RECT 403.150 3.670 407.830 4.280 ;
        RECT 408.670 3.670 413.350 4.280 ;
        RECT 414.190 3.670 418.870 4.280 ;
        RECT 419.710 3.670 424.390 4.280 ;
        RECT 425.230 3.670 429.910 4.280 ;
        RECT 430.750 3.670 435.430 4.280 ;
        RECT 436.270 3.670 440.950 4.280 ;
        RECT 441.790 3.670 446.470 4.280 ;
        RECT 447.310 3.670 451.990 4.280 ;
        RECT 452.830 3.670 457.510 4.280 ;
        RECT 458.350 3.670 463.030 4.280 ;
        RECT 463.870 3.670 468.550 4.280 ;
        RECT 469.390 3.670 474.070 4.280 ;
        RECT 474.910 3.670 479.590 4.280 ;
        RECT 480.430 3.670 485.110 4.280 ;
        RECT 485.950 3.670 490.630 4.280 ;
        RECT 491.470 3.670 496.150 4.280 ;
        RECT 496.990 3.670 501.670 4.280 ;
        RECT 502.510 3.670 507.190 4.280 ;
        RECT 508.030 3.670 512.710 4.280 ;
        RECT 513.550 3.670 518.230 4.280 ;
        RECT 519.070 3.670 523.750 4.280 ;
        RECT 524.590 3.670 529.270 4.280 ;
        RECT 530.110 3.670 534.790 4.280 ;
        RECT 535.630 3.670 540.310 4.280 ;
        RECT 541.150 3.670 545.830 4.280 ;
        RECT 546.670 3.670 551.350 4.280 ;
        RECT 552.190 3.670 556.870 4.280 ;
        RECT 557.710 3.670 562.390 4.280 ;
        RECT 563.230 3.670 567.910 4.280 ;
        RECT 568.750 3.670 573.430 4.280 ;
        RECT 574.270 3.670 578.950 4.280 ;
        RECT 579.790 3.670 584.470 4.280 ;
        RECT 585.310 3.670 589.990 4.280 ;
        RECT 590.830 3.670 595.510 4.280 ;
        RECT 596.350 3.670 601.030 4.280 ;
        RECT 601.870 3.670 606.550 4.280 ;
        RECT 607.390 3.670 612.070 4.280 ;
        RECT 612.910 3.670 617.590 4.280 ;
        RECT 618.430 3.670 623.110 4.280 ;
        RECT 623.950 3.670 628.630 4.280 ;
        RECT 629.470 3.670 634.150 4.280 ;
        RECT 634.990 3.670 639.670 4.280 ;
        RECT 640.510 3.670 645.190 4.280 ;
        RECT 646.030 3.670 650.710 4.280 ;
        RECT 651.550 3.670 656.230 4.280 ;
        RECT 657.070 3.670 661.750 4.280 ;
        RECT 662.590 3.670 667.270 4.280 ;
        RECT 668.110 3.670 672.790 4.280 ;
        RECT 673.630 3.670 678.310 4.280 ;
        RECT 679.150 3.670 683.830 4.280 ;
        RECT 684.670 3.670 689.350 4.280 ;
        RECT 690.190 3.670 694.870 4.280 ;
        RECT 695.710 3.670 700.390 4.280 ;
        RECT 701.230 3.670 705.910 4.280 ;
        RECT 706.750 3.670 711.430 4.280 ;
        RECT 712.270 3.670 716.950 4.280 ;
        RECT 717.790 3.670 722.470 4.280 ;
        RECT 723.310 3.670 727.990 4.280 ;
        RECT 728.830 3.670 733.510 4.280 ;
        RECT 734.350 3.670 739.030 4.280 ;
        RECT 739.870 3.670 744.550 4.280 ;
        RECT 745.390 3.670 750.070 4.280 ;
        RECT 750.910 3.670 755.590 4.280 ;
        RECT 756.430 3.670 761.110 4.280 ;
        RECT 761.950 3.670 766.630 4.280 ;
        RECT 767.470 3.670 772.150 4.280 ;
        RECT 772.990 3.670 777.670 4.280 ;
        RECT 778.510 3.670 783.190 4.280 ;
        RECT 784.030 3.670 788.710 4.280 ;
        RECT 789.550 3.670 794.230 4.280 ;
        RECT 795.070 3.670 799.750 4.280 ;
        RECT 800.590 3.670 805.270 4.280 ;
        RECT 806.110 3.670 810.790 4.280 ;
        RECT 811.630 3.670 816.310 4.280 ;
        RECT 817.150 3.670 821.830 4.280 ;
        RECT 822.670 3.670 827.350 4.280 ;
        RECT 828.190 3.670 832.870 4.280 ;
        RECT 833.710 3.670 838.390 4.280 ;
        RECT 839.230 3.670 843.910 4.280 ;
        RECT 844.750 3.670 849.430 4.280 ;
        RECT 850.270 3.670 854.950 4.280 ;
        RECT 855.790 3.670 860.470 4.280 ;
        RECT 861.310 3.670 865.990 4.280 ;
        RECT 866.830 3.670 871.510 4.280 ;
        RECT 872.350 3.670 877.030 4.280 ;
        RECT 877.870 3.670 882.550 4.280 ;
        RECT 883.390 3.670 888.070 4.280 ;
        RECT 888.910 3.670 893.590 4.280 ;
        RECT 894.430 3.670 899.110 4.280 ;
        RECT 899.950 3.670 904.630 4.280 ;
        RECT 905.470 3.670 910.150 4.280 ;
        RECT 910.990 3.670 915.670 4.280 ;
        RECT 916.510 3.670 921.190 4.280 ;
        RECT 922.030 3.670 926.710 4.280 ;
        RECT 927.550 3.670 932.230 4.280 ;
        RECT 933.070 3.670 937.750 4.280 ;
        RECT 938.590 3.670 943.270 4.280 ;
        RECT 944.110 3.670 948.790 4.280 ;
        RECT 949.630 3.670 954.310 4.280 ;
        RECT 955.150 3.670 959.830 4.280 ;
        RECT 960.670 3.670 965.350 4.280 ;
        RECT 966.190 3.670 970.870 4.280 ;
        RECT 971.710 3.670 976.390 4.280 ;
        RECT 977.230 3.670 981.910 4.280 ;
        RECT 982.750 3.670 987.430 4.280 ;
        RECT 988.270 3.670 992.950 4.280 ;
        RECT 993.790 3.670 998.470 4.280 ;
        RECT 999.310 3.670 1003.990 4.280 ;
        RECT 1004.830 3.670 1009.510 4.280 ;
        RECT 1010.350 3.670 1015.030 4.280 ;
        RECT 1015.870 3.670 1020.550 4.280 ;
        RECT 1021.390 3.670 1026.070 4.280 ;
        RECT 1026.910 3.670 1031.590 4.280 ;
        RECT 1032.430 3.670 1037.110 4.280 ;
        RECT 1037.950 3.670 1042.630 4.280 ;
        RECT 1043.470 3.670 1048.150 4.280 ;
        RECT 1048.990 3.670 1053.670 4.280 ;
        RECT 1054.510 3.670 1059.190 4.280 ;
        RECT 1060.030 3.670 1064.710 4.280 ;
        RECT 1065.550 3.670 1070.230 4.280 ;
        RECT 1071.070 3.670 1075.750 4.280 ;
        RECT 1076.590 3.670 1081.270 4.280 ;
        RECT 1082.110 3.670 1086.790 4.280 ;
        RECT 1087.630 3.670 1092.310 4.280 ;
        RECT 1093.150 3.670 1097.830 4.280 ;
        RECT 1098.670 3.670 1103.350 4.280 ;
        RECT 1104.190 3.670 1108.870 4.280 ;
        RECT 1109.710 3.670 1114.390 4.280 ;
        RECT 1115.230 3.670 1119.910 4.280 ;
        RECT 1120.750 3.670 1125.430 4.280 ;
        RECT 1126.270 3.670 1130.950 4.280 ;
        RECT 1131.790 3.670 1136.470 4.280 ;
        RECT 1137.310 3.670 1141.990 4.280 ;
        RECT 1142.830 3.670 1147.510 4.280 ;
        RECT 1148.350 3.670 1153.030 4.280 ;
        RECT 1153.870 3.670 1158.550 4.280 ;
        RECT 1159.390 3.670 1164.070 4.280 ;
        RECT 1164.910 3.670 1169.590 4.280 ;
        RECT 1170.430 3.670 1175.110 4.280 ;
        RECT 1175.950 3.670 1180.630 4.280 ;
        RECT 1181.470 3.670 1186.150 4.280 ;
        RECT 1186.990 3.670 1191.670 4.280 ;
        RECT 1192.510 3.670 1197.190 4.280 ;
        RECT 1198.030 3.670 1202.710 4.280 ;
        RECT 1203.550 3.670 1208.230 4.280 ;
        RECT 1209.070 3.670 1213.750 4.280 ;
        RECT 1214.590 3.670 1219.270 4.280 ;
        RECT 1220.110 3.670 1224.790 4.280 ;
        RECT 1225.630 3.670 1230.310 4.280 ;
        RECT 1231.150 3.670 1235.830 4.280 ;
        RECT 1236.670 3.670 1241.350 4.280 ;
        RECT 1242.190 3.670 1246.870 4.280 ;
        RECT 1247.710 3.670 1252.390 4.280 ;
        RECT 1253.230 3.670 1257.910 4.280 ;
        RECT 1258.750 3.670 1263.430 4.280 ;
        RECT 1264.270 3.670 1268.950 4.280 ;
        RECT 1269.790 3.670 1274.470 4.280 ;
        RECT 1275.310 3.670 1279.990 4.280 ;
        RECT 1280.830 3.670 1285.510 4.280 ;
        RECT 1286.350 3.670 1291.030 4.280 ;
        RECT 1291.870 3.670 1296.550 4.280 ;
        RECT 1297.390 3.670 1302.070 4.280 ;
        RECT 1302.910 3.670 1307.590 4.280 ;
        RECT 1308.430 3.670 1313.110 4.280 ;
        RECT 1313.950 3.670 1318.630 4.280 ;
        RECT 1319.470 3.670 1324.150 4.280 ;
        RECT 1324.990 3.670 1329.670 4.280 ;
        RECT 1330.510 3.670 1335.190 4.280 ;
        RECT 1336.030 3.670 1340.710 4.280 ;
        RECT 1341.550 3.670 1346.230 4.280 ;
        RECT 1347.070 3.670 1351.750 4.280 ;
        RECT 1352.590 3.670 1357.270 4.280 ;
        RECT 1358.110 3.670 1362.790 4.280 ;
        RECT 1363.630 3.670 1368.310 4.280 ;
        RECT 1369.150 3.670 1373.830 4.280 ;
        RECT 1374.670 3.670 1379.350 4.280 ;
        RECT 1380.190 3.670 1384.870 4.280 ;
        RECT 1385.710 3.670 1390.390 4.280 ;
        RECT 1391.230 3.670 1395.910 4.280 ;
        RECT 1396.750 3.670 1401.430 4.280 ;
        RECT 1402.270 3.670 1406.950 4.280 ;
        RECT 1407.790 3.670 1412.470 4.280 ;
        RECT 1413.310 3.670 1417.990 4.280 ;
        RECT 1418.830 3.670 1423.510 4.280 ;
        RECT 1424.350 3.670 1429.030 4.280 ;
        RECT 1429.870 3.670 1434.550 4.280 ;
        RECT 1435.390 3.670 1440.070 4.280 ;
        RECT 1440.910 3.670 1445.590 4.280 ;
        RECT 1446.430 3.670 1451.110 4.280 ;
        RECT 1451.950 3.670 1456.630 4.280 ;
        RECT 1457.470 3.670 1462.150 4.280 ;
        RECT 1462.990 3.670 1467.670 4.280 ;
        RECT 1468.510 3.670 1473.190 4.280 ;
        RECT 1474.030 3.670 1478.710 4.280 ;
        RECT 1479.550 3.670 1484.230 4.280 ;
        RECT 1485.070 3.670 1489.750 4.280 ;
        RECT 1490.590 3.670 1495.270 4.280 ;
        RECT 1496.110 3.670 1500.790 4.280 ;
        RECT 1501.630 3.670 1506.310 4.280 ;
        RECT 1507.150 3.670 1511.830 4.280 ;
        RECT 1512.670 3.670 1517.350 4.280 ;
        RECT 1518.190 3.670 1522.870 4.280 ;
        RECT 1523.710 3.670 1528.390 4.280 ;
        RECT 1529.230 3.670 1533.910 4.280 ;
        RECT 1534.750 3.670 1539.430 4.280 ;
        RECT 1540.270 3.670 1544.950 4.280 ;
        RECT 1545.790 3.670 1550.470 4.280 ;
        RECT 1551.310 3.670 1555.990 4.280 ;
        RECT 1556.830 3.670 1561.510 4.280 ;
        RECT 1562.350 3.670 1567.030 4.280 ;
        RECT 1567.870 3.670 1572.550 4.280 ;
        RECT 1573.390 3.670 1578.070 4.280 ;
        RECT 1578.910 3.670 1583.590 4.280 ;
        RECT 1584.430 3.670 1589.110 4.280 ;
        RECT 1589.950 3.670 1594.630 4.280 ;
        RECT 1595.470 3.670 1600.150 4.280 ;
        RECT 1600.990 3.670 1605.670 4.280 ;
        RECT 1606.510 3.670 1611.190 4.280 ;
        RECT 1612.030 3.670 1616.710 4.280 ;
        RECT 1617.550 3.670 1622.230 4.280 ;
        RECT 1623.070 3.670 1627.750 4.280 ;
        RECT 1628.590 3.670 1633.270 4.280 ;
        RECT 1634.110 3.670 1638.790 4.280 ;
        RECT 1639.630 3.670 1644.310 4.280 ;
        RECT 1645.150 3.670 1649.830 4.280 ;
        RECT 1650.670 3.670 1655.350 4.280 ;
        RECT 1656.190 3.670 1660.870 4.280 ;
        RECT 1661.710 3.670 1666.390 4.280 ;
        RECT 1667.230 3.670 1671.910 4.280 ;
        RECT 1672.750 3.670 1677.430 4.280 ;
        RECT 1678.270 3.670 1682.950 4.280 ;
        RECT 1683.790 3.670 1688.470 4.280 ;
        RECT 1689.310 3.670 1693.990 4.280 ;
        RECT 1694.830 3.670 1699.510 4.280 ;
        RECT 1700.350 3.670 1705.030 4.280 ;
        RECT 1705.870 3.670 1710.550 4.280 ;
        RECT 1711.390 3.670 1716.070 4.280 ;
        RECT 1716.910 3.670 1721.590 4.280 ;
        RECT 1722.430 3.670 1727.110 4.280 ;
        RECT 1727.950 3.670 1732.630 4.280 ;
        RECT 1733.470 3.670 1738.150 4.280 ;
        RECT 1738.990 3.670 1743.670 4.280 ;
        RECT 1744.510 3.670 1749.190 4.280 ;
        RECT 1750.030 3.670 1754.710 4.280 ;
        RECT 1755.550 3.670 1760.230 4.280 ;
        RECT 1761.070 3.670 1765.750 4.280 ;
        RECT 1766.590 3.670 1771.270 4.280 ;
        RECT 1772.110 3.670 1776.790 4.280 ;
        RECT 1777.630 3.670 1782.310 4.280 ;
        RECT 1783.150 3.670 1787.830 4.280 ;
        RECT 1788.670 3.670 1793.350 4.280 ;
        RECT 1794.190 3.670 1798.870 4.280 ;
        RECT 1799.710 3.670 1804.390 4.280 ;
        RECT 1805.230 3.670 1809.910 4.280 ;
        RECT 1810.750 3.670 1815.430 4.280 ;
        RECT 1816.270 3.670 1820.950 4.280 ;
        RECT 1821.790 3.670 1826.470 4.280 ;
        RECT 1827.310 3.670 1831.990 4.280 ;
        RECT 1832.830 3.670 1837.510 4.280 ;
        RECT 1838.350 3.670 1843.030 4.280 ;
        RECT 1843.870 3.670 1848.550 4.280 ;
        RECT 1849.390 3.670 1854.070 4.280 ;
        RECT 1854.910 3.670 1859.590 4.280 ;
        RECT 1860.430 3.670 1865.110 4.280 ;
        RECT 1865.950 3.670 1870.630 4.280 ;
        RECT 1871.470 3.670 1876.150 4.280 ;
        RECT 1876.990 3.670 1881.670 4.280 ;
        RECT 1882.510 3.670 1887.190 4.280 ;
        RECT 1888.030 3.670 1892.710 4.280 ;
        RECT 1893.550 3.670 1898.230 4.280 ;
        RECT 1899.070 3.670 1903.750 4.280 ;
        RECT 1904.590 3.670 1909.270 4.280 ;
        RECT 1910.110 3.670 1914.790 4.280 ;
        RECT 1915.630 3.670 1920.310 4.280 ;
        RECT 1921.150 3.670 1925.830 4.280 ;
        RECT 1926.670 3.670 1931.350 4.280 ;
        RECT 1932.190 3.670 1936.870 4.280 ;
        RECT 1937.710 3.670 1942.390 4.280 ;
        RECT 1943.230 3.670 1947.910 4.280 ;
        RECT 1948.750 3.670 1953.430 4.280 ;
        RECT 1954.270 3.670 1958.950 4.280 ;
        RECT 1959.790 3.670 1964.470 4.280 ;
        RECT 1965.310 3.670 1969.990 4.280 ;
        RECT 1970.830 3.670 1975.510 4.280 ;
        RECT 1976.350 3.670 1981.030 4.280 ;
        RECT 1981.870 3.670 1986.550 4.280 ;
        RECT 1987.390 3.670 1992.070 4.280 ;
        RECT 1992.910 3.670 1997.590 4.280 ;
        RECT 1998.430 3.670 2003.110 4.280 ;
        RECT 2003.950 3.670 2008.630 4.280 ;
        RECT 2009.470 3.670 2014.150 4.280 ;
        RECT 2014.990 3.670 2019.670 4.280 ;
        RECT 2020.510 3.670 2025.190 4.280 ;
        RECT 2026.030 3.670 2030.710 4.280 ;
        RECT 2031.550 3.670 2036.230 4.280 ;
        RECT 2037.070 3.670 2041.750 4.280 ;
        RECT 2042.590 3.670 2047.270 4.280 ;
        RECT 2048.110 3.670 2052.790 4.280 ;
        RECT 2053.630 3.670 2058.310 4.280 ;
        RECT 2059.150 3.670 2063.830 4.280 ;
        RECT 2064.670 3.670 2069.350 4.280 ;
        RECT 2070.190 3.670 2074.870 4.280 ;
        RECT 2075.710 3.670 2080.390 4.280 ;
        RECT 2081.230 3.670 2085.910 4.280 ;
        RECT 2086.750 3.670 2091.430 4.280 ;
        RECT 2092.270 3.670 2096.950 4.280 ;
        RECT 2097.790 3.670 2102.470 4.280 ;
        RECT 2103.310 3.670 2107.990 4.280 ;
        RECT 2108.830 3.670 2113.510 4.280 ;
        RECT 2114.350 3.670 2119.030 4.280 ;
        RECT 2119.870 3.670 2124.550 4.280 ;
        RECT 2125.390 3.670 2130.070 4.280 ;
        RECT 2130.910 3.670 2135.590 4.280 ;
        RECT 2136.430 3.670 2141.110 4.280 ;
        RECT 2141.950 3.670 2146.630 4.280 ;
        RECT 2147.470 3.670 2152.150 4.280 ;
        RECT 2152.990 3.670 2157.670 4.280 ;
        RECT 2158.510 3.670 2163.190 4.280 ;
        RECT 2164.030 3.670 2168.710 4.280 ;
        RECT 2169.550 3.670 2174.230 4.280 ;
        RECT 2175.070 3.670 2179.750 4.280 ;
        RECT 2180.590 3.670 2185.270 4.280 ;
        RECT 2186.110 3.670 2190.790 4.280 ;
        RECT 2191.630 3.670 2196.310 4.280 ;
        RECT 2197.150 3.670 2201.830 4.280 ;
        RECT 2202.670 3.670 2207.350 4.280 ;
        RECT 2208.190 3.670 2212.870 4.280 ;
        RECT 2213.710 3.670 2218.390 4.280 ;
        RECT 2219.230 3.670 2223.910 4.280 ;
        RECT 2224.750 3.670 2229.430 4.280 ;
        RECT 2230.270 3.670 2234.950 4.280 ;
        RECT 2235.790 3.670 2240.470 4.280 ;
        RECT 2241.310 3.670 2245.990 4.280 ;
        RECT 2246.830 3.670 2251.510 4.280 ;
        RECT 2252.350 3.670 2257.030 4.280 ;
        RECT 2257.870 3.670 2262.550 4.280 ;
        RECT 2263.390 3.670 2268.070 4.280 ;
        RECT 2268.910 3.670 2273.590 4.280 ;
        RECT 2274.430 3.670 2279.110 4.280 ;
        RECT 2279.950 3.670 2284.630 4.280 ;
        RECT 2285.470 3.670 2290.150 4.280 ;
        RECT 2290.990 3.670 2295.670 4.280 ;
        RECT 2296.510 3.670 2301.190 4.280 ;
        RECT 2302.030 3.670 2306.710 4.280 ;
        RECT 2307.550 3.670 2312.230 4.280 ;
        RECT 2313.070 3.670 2317.750 4.280 ;
        RECT 2318.590 3.670 2323.270 4.280 ;
        RECT 2324.110 3.670 2328.790 4.280 ;
        RECT 2329.630 3.670 2334.310 4.280 ;
        RECT 2335.150 3.670 2339.830 4.280 ;
        RECT 2340.670 3.670 2345.350 4.280 ;
        RECT 2346.190 3.670 2350.870 4.280 ;
        RECT 2351.710 3.670 2356.390 4.280 ;
        RECT 2357.230 3.670 2361.910 4.280 ;
        RECT 2362.750 3.670 2367.430 4.280 ;
        RECT 2368.270 3.670 2372.950 4.280 ;
        RECT 2373.790 3.670 2378.470 4.280 ;
        RECT 2379.310 3.670 2383.990 4.280 ;
        RECT 2384.830 3.670 2389.510 4.280 ;
        RECT 2390.350 3.670 2395.030 4.280 ;
        RECT 2395.870 3.670 2400.550 4.280 ;
        RECT 2401.390 3.670 2406.070 4.280 ;
        RECT 2406.910 3.670 2411.590 4.280 ;
        RECT 2412.430 3.670 2417.110 4.280 ;
        RECT 2417.950 3.670 2422.630 4.280 ;
        RECT 2423.470 3.670 2428.150 4.280 ;
        RECT 2428.990 3.670 2433.670 4.280 ;
        RECT 2434.510 3.670 2439.190 4.280 ;
        RECT 2440.030 3.670 2444.710 4.280 ;
        RECT 2445.550 3.670 2450.230 4.280 ;
        RECT 2451.070 3.670 2455.750 4.280 ;
        RECT 2456.590 3.670 2461.270 4.280 ;
        RECT 2462.110 3.670 2466.790 4.280 ;
        RECT 2467.630 3.670 2472.310 4.280 ;
        RECT 2473.150 3.670 2477.830 4.280 ;
        RECT 2478.670 3.670 2483.350 4.280 ;
        RECT 2484.190 3.670 2488.870 4.280 ;
        RECT 2489.710 3.670 2494.390 4.280 ;
        RECT 2495.230 3.670 2499.910 4.280 ;
        RECT 2500.750 3.670 2505.430 4.280 ;
        RECT 2506.270 3.670 2510.950 4.280 ;
        RECT 2511.790 3.670 2516.470 4.280 ;
        RECT 2517.310 3.670 2521.990 4.280 ;
        RECT 2522.830 3.670 2527.510 4.280 ;
        RECT 2528.350 3.670 2533.030 4.280 ;
        RECT 2533.870 3.670 2538.550 4.280 ;
        RECT 2539.390 3.670 2544.070 4.280 ;
        RECT 2544.910 3.670 2549.590 4.280 ;
        RECT 2550.430 3.670 2555.110 4.280 ;
        RECT 2555.950 3.670 2560.630 4.280 ;
        RECT 2561.470 3.670 2566.150 4.280 ;
        RECT 2566.990 3.670 2571.670 4.280 ;
        RECT 2572.510 3.670 2577.190 4.280 ;
        RECT 2578.030 3.670 2582.710 4.280 ;
        RECT 2583.550 3.670 2588.230 4.280 ;
        RECT 2589.070 3.670 2593.750 4.280 ;
        RECT 2594.590 3.670 2599.270 4.280 ;
        RECT 2600.110 3.670 2604.790 4.280 ;
        RECT 2605.630 3.670 2610.310 4.280 ;
        RECT 2611.150 3.670 2615.830 4.280 ;
        RECT 2616.670 3.670 2621.350 4.280 ;
        RECT 2622.190 3.670 2626.870 4.280 ;
        RECT 2627.710 3.670 2632.390 4.280 ;
        RECT 2633.230 3.670 2637.910 4.280 ;
        RECT 2638.750 3.670 2643.430 4.280 ;
        RECT 2644.270 3.670 2648.950 4.280 ;
        RECT 2649.790 3.670 2654.470 4.280 ;
        RECT 2655.310 3.670 2659.990 4.280 ;
        RECT 2660.830 3.670 2665.510 4.280 ;
        RECT 2666.350 3.670 2671.030 4.280 ;
        RECT 2671.870 3.670 2676.550 4.280 ;
        RECT 2677.390 3.670 2682.070 4.280 ;
        RECT 2682.910 3.670 2687.590 4.280 ;
        RECT 2688.430 3.670 2693.110 4.280 ;
        RECT 2693.950 3.670 2698.630 4.280 ;
        RECT 2699.470 3.670 2704.150 4.280 ;
        RECT 2704.990 3.670 2709.670 4.280 ;
        RECT 2710.510 3.670 2715.190 4.280 ;
        RECT 2716.030 3.670 2720.710 4.280 ;
        RECT 2721.550 3.670 2726.230 4.280 ;
        RECT 2727.070 3.670 2731.750 4.280 ;
        RECT 2732.590 3.670 2737.270 4.280 ;
        RECT 2738.110 3.670 2742.790 4.280 ;
        RECT 2743.630 3.670 2748.310 4.280 ;
        RECT 2749.150 3.670 2753.830 4.280 ;
        RECT 2754.670 3.670 2759.350 4.280 ;
        RECT 2760.190 3.670 2764.870 4.280 ;
        RECT 2765.710 3.670 2770.390 4.280 ;
        RECT 2771.230 3.670 2775.910 4.280 ;
        RECT 2776.750 3.670 2781.430 4.280 ;
        RECT 2782.270 3.670 2786.950 4.280 ;
        RECT 2787.790 3.670 2853.740 4.280 ;
      LAYER met3 ;
        RECT 1.905 3396.960 2853.315 3421.925 ;
        RECT 1.905 3395.560 2849.625 3396.960 ;
        RECT 1.905 3392.880 2853.315 3395.560 ;
        RECT 4.400 3391.480 2853.315 3392.880 ;
        RECT 1.905 3332.360 2853.315 3391.480 ;
        RECT 1.905 3330.960 2849.625 3332.360 ;
        RECT 1.905 3329.640 2853.315 3330.960 ;
        RECT 4.400 3328.240 2853.315 3329.640 ;
        RECT 1.905 3267.760 2853.315 3328.240 ;
        RECT 1.905 3266.400 2849.625 3267.760 ;
        RECT 4.400 3266.360 2849.625 3266.400 ;
        RECT 4.400 3265.000 2853.315 3266.360 ;
        RECT 1.905 3203.160 2853.315 3265.000 ;
        RECT 4.400 3201.760 2849.625 3203.160 ;
        RECT 1.905 3139.920 2853.315 3201.760 ;
        RECT 4.400 3138.560 2853.315 3139.920 ;
        RECT 4.400 3138.520 2849.625 3138.560 ;
        RECT 1.905 3137.160 2849.625 3138.520 ;
        RECT 1.905 3076.680 2853.315 3137.160 ;
        RECT 4.400 3075.280 2853.315 3076.680 ;
        RECT 1.905 3073.960 2853.315 3075.280 ;
        RECT 1.905 3072.560 2849.625 3073.960 ;
        RECT 1.905 3013.440 2853.315 3072.560 ;
        RECT 4.400 3012.040 2853.315 3013.440 ;
        RECT 1.905 3009.360 2853.315 3012.040 ;
        RECT 1.905 3007.960 2849.625 3009.360 ;
        RECT 1.905 2950.200 2853.315 3007.960 ;
        RECT 4.400 2948.800 2853.315 2950.200 ;
        RECT 1.905 2944.760 2853.315 2948.800 ;
        RECT 1.905 2943.360 2849.625 2944.760 ;
        RECT 1.905 2886.960 2853.315 2943.360 ;
        RECT 4.400 2885.560 2853.315 2886.960 ;
        RECT 1.905 2880.160 2853.315 2885.560 ;
        RECT 1.905 2878.760 2849.625 2880.160 ;
        RECT 1.905 2823.720 2853.315 2878.760 ;
        RECT 4.400 2822.320 2853.315 2823.720 ;
        RECT 1.905 2815.560 2853.315 2822.320 ;
        RECT 1.905 2814.160 2849.625 2815.560 ;
        RECT 1.905 2760.480 2853.315 2814.160 ;
        RECT 4.400 2759.080 2853.315 2760.480 ;
        RECT 1.905 2750.960 2853.315 2759.080 ;
        RECT 1.905 2749.560 2849.625 2750.960 ;
        RECT 1.905 2697.240 2853.315 2749.560 ;
        RECT 4.400 2695.840 2853.315 2697.240 ;
        RECT 1.905 2686.360 2853.315 2695.840 ;
        RECT 1.905 2684.960 2849.625 2686.360 ;
        RECT 1.905 2634.000 2853.315 2684.960 ;
        RECT 4.400 2632.600 2853.315 2634.000 ;
        RECT 1.905 2621.760 2853.315 2632.600 ;
        RECT 1.905 2620.360 2849.625 2621.760 ;
        RECT 1.905 2570.760 2853.315 2620.360 ;
        RECT 4.400 2569.360 2853.315 2570.760 ;
        RECT 1.905 2557.160 2853.315 2569.360 ;
        RECT 1.905 2555.760 2849.625 2557.160 ;
        RECT 1.905 2507.520 2853.315 2555.760 ;
        RECT 4.400 2506.120 2853.315 2507.520 ;
        RECT 1.905 2492.560 2853.315 2506.120 ;
        RECT 1.905 2491.160 2849.625 2492.560 ;
        RECT 1.905 2444.280 2853.315 2491.160 ;
        RECT 4.400 2442.880 2853.315 2444.280 ;
        RECT 1.905 2427.960 2853.315 2442.880 ;
        RECT 1.905 2426.560 2849.625 2427.960 ;
        RECT 1.905 2381.040 2853.315 2426.560 ;
        RECT 4.400 2379.640 2853.315 2381.040 ;
        RECT 1.905 2363.360 2853.315 2379.640 ;
        RECT 1.905 2361.960 2849.625 2363.360 ;
        RECT 1.905 2317.800 2853.315 2361.960 ;
        RECT 4.400 2316.400 2853.315 2317.800 ;
        RECT 1.905 2298.760 2853.315 2316.400 ;
        RECT 1.905 2297.360 2849.625 2298.760 ;
        RECT 1.905 2254.560 2853.315 2297.360 ;
        RECT 4.400 2253.160 2853.315 2254.560 ;
        RECT 1.905 2234.160 2853.315 2253.160 ;
        RECT 1.905 2232.760 2849.625 2234.160 ;
        RECT 1.905 2191.320 2853.315 2232.760 ;
        RECT 4.400 2189.920 2853.315 2191.320 ;
        RECT 1.905 2169.560 2853.315 2189.920 ;
        RECT 1.905 2168.160 2849.625 2169.560 ;
        RECT 1.905 2128.080 2853.315 2168.160 ;
        RECT 4.400 2126.680 2853.315 2128.080 ;
        RECT 1.905 2104.960 2853.315 2126.680 ;
        RECT 1.905 2103.560 2849.625 2104.960 ;
        RECT 1.905 2064.840 2853.315 2103.560 ;
        RECT 4.400 2063.440 2853.315 2064.840 ;
        RECT 1.905 2040.360 2853.315 2063.440 ;
        RECT 1.905 2038.960 2849.625 2040.360 ;
        RECT 1.905 2001.600 2853.315 2038.960 ;
        RECT 4.400 2000.200 2853.315 2001.600 ;
        RECT 1.905 1975.760 2853.315 2000.200 ;
        RECT 1.905 1974.360 2849.625 1975.760 ;
        RECT 1.905 1938.360 2853.315 1974.360 ;
        RECT 4.400 1936.960 2853.315 1938.360 ;
        RECT 1.905 1911.160 2853.315 1936.960 ;
        RECT 1.905 1909.760 2849.625 1911.160 ;
        RECT 1.905 1875.120 2853.315 1909.760 ;
        RECT 4.400 1873.720 2853.315 1875.120 ;
        RECT 1.905 1846.560 2853.315 1873.720 ;
        RECT 1.905 1845.160 2849.625 1846.560 ;
        RECT 1.905 1811.880 2853.315 1845.160 ;
        RECT 4.400 1810.480 2853.315 1811.880 ;
        RECT 1.905 1781.960 2853.315 1810.480 ;
        RECT 1.905 1780.560 2849.625 1781.960 ;
        RECT 1.905 1748.640 2853.315 1780.560 ;
        RECT 4.400 1747.240 2853.315 1748.640 ;
        RECT 1.905 1717.360 2853.315 1747.240 ;
        RECT 1.905 1715.960 2849.625 1717.360 ;
        RECT 1.905 1685.400 2853.315 1715.960 ;
        RECT 4.400 1684.000 2853.315 1685.400 ;
        RECT 1.905 1652.760 2853.315 1684.000 ;
        RECT 1.905 1651.360 2849.625 1652.760 ;
        RECT 1.905 1622.160 2853.315 1651.360 ;
        RECT 4.400 1620.760 2853.315 1622.160 ;
        RECT 1.905 1588.160 2853.315 1620.760 ;
        RECT 1.905 1586.760 2849.625 1588.160 ;
        RECT 1.905 1558.920 2853.315 1586.760 ;
        RECT 4.400 1557.520 2853.315 1558.920 ;
        RECT 1.905 1523.560 2853.315 1557.520 ;
        RECT 1.905 1522.160 2849.625 1523.560 ;
        RECT 1.905 1495.680 2853.315 1522.160 ;
        RECT 4.400 1494.280 2853.315 1495.680 ;
        RECT 1.905 1458.960 2853.315 1494.280 ;
        RECT 1.905 1457.560 2849.625 1458.960 ;
        RECT 1.905 1432.440 2853.315 1457.560 ;
        RECT 4.400 1431.040 2853.315 1432.440 ;
        RECT 1.905 1394.360 2853.315 1431.040 ;
        RECT 1.905 1392.960 2849.625 1394.360 ;
        RECT 1.905 1369.200 2853.315 1392.960 ;
        RECT 4.400 1367.800 2853.315 1369.200 ;
        RECT 1.905 1329.760 2853.315 1367.800 ;
        RECT 1.905 1328.360 2849.625 1329.760 ;
        RECT 1.905 1305.960 2853.315 1328.360 ;
        RECT 4.400 1304.560 2853.315 1305.960 ;
        RECT 1.905 1265.160 2853.315 1304.560 ;
        RECT 1.905 1263.760 2849.625 1265.160 ;
        RECT 1.905 1242.720 2853.315 1263.760 ;
        RECT 4.400 1241.320 2853.315 1242.720 ;
        RECT 1.905 1200.560 2853.315 1241.320 ;
        RECT 1.905 1199.160 2849.625 1200.560 ;
        RECT 1.905 1179.480 2853.315 1199.160 ;
        RECT 4.400 1178.080 2853.315 1179.480 ;
        RECT 1.905 1135.960 2853.315 1178.080 ;
        RECT 1.905 1134.560 2849.625 1135.960 ;
        RECT 1.905 1116.240 2853.315 1134.560 ;
        RECT 4.400 1114.840 2853.315 1116.240 ;
        RECT 1.905 1071.360 2853.315 1114.840 ;
        RECT 1.905 1069.960 2849.625 1071.360 ;
        RECT 1.905 1053.000 2853.315 1069.960 ;
        RECT 4.400 1051.600 2853.315 1053.000 ;
        RECT 1.905 1006.760 2853.315 1051.600 ;
        RECT 1.905 1005.360 2849.625 1006.760 ;
        RECT 1.905 989.760 2853.315 1005.360 ;
        RECT 4.400 988.360 2853.315 989.760 ;
        RECT 1.905 942.160 2853.315 988.360 ;
        RECT 1.905 940.760 2849.625 942.160 ;
        RECT 1.905 926.520 2853.315 940.760 ;
        RECT 4.400 925.120 2853.315 926.520 ;
        RECT 1.905 877.560 2853.315 925.120 ;
        RECT 1.905 876.160 2849.625 877.560 ;
        RECT 1.905 863.280 2853.315 876.160 ;
        RECT 4.400 861.880 2853.315 863.280 ;
        RECT 1.905 812.960 2853.315 861.880 ;
        RECT 1.905 811.560 2849.625 812.960 ;
        RECT 1.905 800.040 2853.315 811.560 ;
        RECT 4.400 798.640 2853.315 800.040 ;
        RECT 1.905 748.360 2853.315 798.640 ;
        RECT 1.905 746.960 2849.625 748.360 ;
        RECT 1.905 736.800 2853.315 746.960 ;
        RECT 4.400 735.400 2853.315 736.800 ;
        RECT 1.905 683.760 2853.315 735.400 ;
        RECT 1.905 682.360 2849.625 683.760 ;
        RECT 1.905 673.560 2853.315 682.360 ;
        RECT 4.400 672.160 2853.315 673.560 ;
        RECT 1.905 619.160 2853.315 672.160 ;
        RECT 1.905 617.760 2849.625 619.160 ;
        RECT 1.905 610.320 2853.315 617.760 ;
        RECT 4.400 608.920 2853.315 610.320 ;
        RECT 1.905 554.560 2853.315 608.920 ;
        RECT 1.905 553.160 2849.625 554.560 ;
        RECT 1.905 547.080 2853.315 553.160 ;
        RECT 4.400 545.680 2853.315 547.080 ;
        RECT 1.905 489.960 2853.315 545.680 ;
        RECT 1.905 488.560 2849.625 489.960 ;
        RECT 1.905 483.840 2853.315 488.560 ;
        RECT 4.400 482.440 2853.315 483.840 ;
        RECT 1.905 425.360 2853.315 482.440 ;
        RECT 1.905 423.960 2849.625 425.360 ;
        RECT 1.905 420.600 2853.315 423.960 ;
        RECT 4.400 419.200 2853.315 420.600 ;
        RECT 1.905 360.760 2853.315 419.200 ;
        RECT 1.905 359.360 2849.625 360.760 ;
        RECT 1.905 357.360 2853.315 359.360 ;
        RECT 4.400 355.960 2853.315 357.360 ;
        RECT 1.905 296.160 2853.315 355.960 ;
        RECT 1.905 294.760 2849.625 296.160 ;
        RECT 1.905 294.120 2853.315 294.760 ;
        RECT 4.400 292.720 2853.315 294.120 ;
        RECT 1.905 231.560 2853.315 292.720 ;
        RECT 1.905 230.880 2849.625 231.560 ;
        RECT 4.400 230.160 2849.625 230.880 ;
        RECT 4.400 229.480 2853.315 230.160 ;
        RECT 1.905 167.640 2853.315 229.480 ;
        RECT 4.400 166.960 2853.315 167.640 ;
        RECT 4.400 166.240 2849.625 166.960 ;
        RECT 1.905 165.560 2849.625 166.240 ;
        RECT 1.905 104.400 2853.315 165.560 ;
        RECT 4.400 103.000 2853.315 104.400 ;
        RECT 1.905 102.360 2853.315 103.000 ;
        RECT 1.905 100.960 2849.625 102.360 ;
        RECT 1.905 41.160 2853.315 100.960 ;
        RECT 4.400 39.760 2853.315 41.160 ;
        RECT 1.905 37.760 2853.315 39.760 ;
        RECT 1.905 36.360 2849.625 37.760 ;
        RECT 1.905 10.715 2853.315 36.360 ;
      LAYER met4 ;
        RECT 2.135 17.175 20.640 3420.225 ;
        RECT 23.040 17.175 97.440 3420.225 ;
        RECT 99.840 17.175 174.240 3420.225 ;
        RECT 176.640 17.175 251.040 3420.225 ;
        RECT 253.440 17.175 327.840 3420.225 ;
        RECT 330.240 17.175 404.640 3420.225 ;
        RECT 407.040 17.175 481.440 3420.225 ;
        RECT 483.840 17.175 558.240 3420.225 ;
        RECT 560.640 17.175 635.040 3420.225 ;
        RECT 637.440 17.175 711.840 3420.225 ;
        RECT 714.240 17.175 788.640 3420.225 ;
        RECT 791.040 17.175 865.440 3420.225 ;
        RECT 867.840 17.175 942.240 3420.225 ;
        RECT 944.640 17.175 1019.040 3420.225 ;
        RECT 1021.440 17.175 1095.840 3420.225 ;
        RECT 1098.240 17.175 1172.640 3420.225 ;
        RECT 1175.040 17.175 1249.440 3420.225 ;
        RECT 1251.840 17.175 1326.240 3420.225 ;
        RECT 1328.640 17.175 1403.040 3420.225 ;
        RECT 1405.440 17.175 1479.840 3420.225 ;
        RECT 1482.240 17.175 1556.640 3420.225 ;
        RECT 1559.040 17.175 1633.440 3420.225 ;
        RECT 1635.840 17.175 1710.240 3420.225 ;
        RECT 1712.640 17.175 1787.040 3420.225 ;
        RECT 1789.440 17.175 1863.840 3420.225 ;
        RECT 1866.240 17.175 1940.640 3420.225 ;
        RECT 1943.040 17.175 2017.440 3420.225 ;
        RECT 2019.840 17.175 2094.240 3420.225 ;
        RECT 2096.640 17.175 2171.040 3420.225 ;
        RECT 2173.440 17.175 2247.840 3420.225 ;
        RECT 2250.240 17.175 2324.640 3420.225 ;
        RECT 2327.040 17.175 2401.440 3420.225 ;
        RECT 2403.840 17.175 2478.240 3420.225 ;
        RECT 2480.640 17.175 2555.040 3420.225 ;
        RECT 2557.440 17.175 2631.840 3420.225 ;
        RECT 2634.240 17.175 2708.640 3420.225 ;
        RECT 2711.040 17.175 2785.440 3420.225 ;
        RECT 2787.840 17.175 2842.505 3420.225 ;
  END
END rift2Wrap
END LIBRARY

