magic
tech sky130A
magscale 1 2
timestamp 1672367698
<< metal1 >>
rect 201494 702992 201500 703044
rect 201552 703032 201558 703044
rect 202782 703032 202788 703044
rect 201552 703004 202788 703032
rect 201552 702992 201558 703004
rect 202782 702992 202788 703004
rect 202840 702992 202846 703044
rect 105446 700884 105452 700936
rect 105504 700924 105510 700936
rect 109034 700924 109040 700936
rect 105504 700896 109040 700924
rect 105504 700884 105510 700896
rect 109034 700884 109040 700896
rect 109092 700884 109098 700936
rect 89162 700680 89168 700732
rect 89220 700720 89226 700732
rect 93026 700720 93032 700732
rect 89220 700692 93032 700720
rect 89220 700680 89226 700692
rect 93026 700680 93032 700692
rect 93084 700680 93090 700732
rect 56778 700476 56784 700528
rect 56836 700516 56842 700528
rect 61378 700516 61384 700528
rect 56836 700488 61384 700516
rect 56836 700476 56842 700488
rect 61378 700476 61384 700488
rect 61436 700476 61442 700528
rect 40494 700340 40500 700392
rect 40552 700380 40558 700392
rect 44174 700380 44180 700392
rect 40552 700352 44180 700380
rect 40552 700340 40558 700352
rect 44174 700340 44180 700352
rect 44232 700340 44238 700392
rect 8110 700272 8116 700324
rect 8168 700312 8174 700324
rect 13906 700312 13912 700324
rect 8168 700284 13912 700312
rect 8168 700272 8174 700284
rect 13906 700272 13912 700284
rect 13964 700272 13970 700324
rect 24302 699660 24308 699712
rect 24360 699700 24366 699712
rect 28258 699700 28264 699712
rect 24360 699672 28264 699700
rect 24360 699660 24366 699672
rect 28258 699660 28264 699672
rect 28316 699660 28322 699712
rect 72970 699660 72976 699712
rect 73028 699700 73034 699712
rect 76098 699700 76104 699712
rect 73028 699672 76104 699700
rect 73028 699660 73034 699672
rect 76098 699660 76104 699672
rect 76156 699660 76162 699712
rect 137830 699660 137836 699712
rect 137888 699700 137894 699712
rect 140774 699700 140780 699712
rect 137888 699672 140780 699700
rect 137888 699660 137894 699672
rect 140774 699660 140780 699672
rect 140832 699660 140838 699712
rect 298738 699660 298744 699712
rect 298796 699700 298802 699712
rect 300118 699700 300124 699712
rect 298796 699672 300124 699700
rect 298796 699660 298802 699672
rect 300118 699660 300124 699672
rect 300176 699660 300182 699712
rect 314654 699660 314660 699712
rect 314712 699700 314718 699712
rect 316310 699700 316316 699712
rect 314712 699672 316316 699700
rect 314712 699660 314718 699672
rect 316310 699660 316316 699672
rect 316368 699660 316374 699712
rect 330386 699660 330392 699712
rect 330444 699700 330450 699712
rect 332502 699700 332508 699712
rect 330444 699672 332508 699700
rect 330444 699660 330450 699672
rect 332502 699660 332508 699672
rect 332560 699660 332566 699712
rect 346394 699660 346400 699712
rect 346452 699700 346458 699712
rect 348786 699700 348792 699712
rect 346452 699672 348792 699700
rect 346452 699660 346458 699672
rect 348786 699660 348792 699672
rect 348844 699660 348850 699712
rect 362034 699660 362040 699712
rect 362092 699700 362098 699712
rect 364978 699700 364984 699712
rect 362092 699672 364984 699700
rect 362092 699660 362098 699672
rect 364978 699660 364984 699672
rect 365036 699660 365042 699712
rect 378134 699660 378140 699712
rect 378192 699700 378198 699712
rect 381170 699700 381176 699712
rect 378192 699672 381176 699700
rect 378192 699660 378198 699672
rect 381170 699660 381176 699672
rect 381228 699660 381234 699712
rect 393682 699660 393688 699712
rect 393740 699700 393746 699712
rect 397454 699700 397460 699712
rect 393740 699672 397460 699700
rect 393740 699660 393746 699672
rect 397454 699660 397460 699672
rect 397512 699660 397518 699712
rect 409874 699660 409880 699712
rect 409932 699700 409938 699712
rect 413646 699700 413652 699712
rect 409932 699672 413652 699700
rect 409932 699660 409938 699672
rect 413646 699660 413652 699672
rect 413704 699660 413710 699712
rect 425330 699660 425336 699712
rect 425388 699700 425394 699712
rect 429838 699700 429844 699712
rect 425388 699672 429844 699700
rect 425388 699660 425394 699672
rect 429838 699660 429844 699672
rect 429896 699660 429902 699712
rect 441614 699660 441620 699712
rect 441672 699700 441678 699712
rect 446122 699700 446128 699712
rect 441672 699672 446128 699700
rect 441672 699660 441678 699672
rect 446122 699660 446128 699672
rect 446180 699660 446186 699712
rect 574094 699660 574100 699712
rect 574152 699700 574158 699712
rect 575842 699700 575848 699712
rect 574152 699672 575848 699700
rect 574152 699660 574158 699672
rect 575842 699660 575848 699672
rect 575900 699660 575906 699712
rect 28258 695444 28264 695496
rect 28316 695484 28322 695496
rect 30190 695484 30196 695496
rect 28316 695456 30196 695484
rect 28316 695444 28322 695456
rect 30190 695444 30196 695456
rect 30248 695444 30254 695496
rect 76098 695444 76104 695496
rect 76156 695484 76162 695496
rect 77662 695484 77668 695496
rect 76156 695456 77668 695484
rect 76156 695444 76162 695456
rect 77662 695444 77668 695456
rect 77720 695444 77726 695496
rect 153194 695444 153200 695496
rect 153252 695484 153258 695496
rect 156782 695484 156788 695496
rect 153252 695456 156788 695484
rect 153252 695444 153258 695456
rect 156782 695444 156788 695456
rect 156840 695444 156846 695496
rect 186498 695444 186504 695496
rect 186556 695484 186562 695496
rect 188430 695484 188436 695496
rect 186556 695456 188436 695484
rect 186556 695444 186562 695456
rect 188430 695444 188436 695456
rect 188488 695444 188494 695496
rect 201494 695444 201500 695496
rect 201552 695484 201558 695496
rect 204254 695484 204260 695496
rect 201552 695456 204260 695484
rect 201552 695444 201558 695456
rect 204254 695444 204260 695456
rect 204312 695444 204318 695496
rect 520734 695444 520740 695496
rect 520792 695484 520798 695496
rect 527174 695484 527180 695496
rect 520792 695456 527180 695484
rect 520792 695444 520798 695456
rect 527174 695444 527180 695456
rect 527232 695444 527238 695496
rect 473262 695376 473268 695428
rect 473320 695416 473326 695428
rect 477494 695416 477500 695428
rect 473320 695388 477500 695416
rect 473320 695376 473326 695388
rect 477494 695376 477500 695388
rect 477552 695376 477558 695428
rect 568206 695240 568212 695292
rect 568264 695280 568270 695292
rect 574094 695280 574100 695292
rect 568264 695252 574100 695280
rect 568264 695240 568270 695252
rect 574094 695240 574100 695252
rect 574152 695240 574158 695292
rect 489086 694764 489092 694816
rect 489144 694804 489150 694816
rect 494054 694804 494060 694816
rect 489144 694776 494060 694804
rect 489144 694764 489150 694776
rect 494054 694764 494060 694776
rect 494112 694764 494118 694816
rect 536558 694764 536564 694816
rect 536616 694804 536622 694816
rect 542354 694804 542360 694816
rect 536616 694776 542360 694804
rect 536616 694764 536622 694776
rect 542354 694764 542360 694776
rect 542412 694764 542418 694816
rect 44174 694152 44180 694204
rect 44232 694192 44238 694204
rect 46014 694192 46020 694204
rect 44232 694164 46020 694192
rect 44232 694152 44238 694164
rect 46014 694152 46020 694164
rect 46072 694152 46078 694204
rect 121638 694152 121644 694204
rect 121696 694192 121702 694204
rect 125134 694192 125140 694204
rect 121696 694164 125140 694192
rect 121696 694152 121702 694164
rect 125134 694152 125140 694164
rect 125192 694152 125198 694204
rect 169754 694152 169760 694204
rect 169812 694192 169818 694204
rect 172606 694192 172612 694204
rect 169812 694164 172612 694192
rect 169812 694152 169818 694164
rect 172606 694152 172612 694164
rect 172664 694152 172670 694204
rect 218054 694152 218060 694204
rect 218112 694192 218118 694204
rect 220078 694192 220084 694204
rect 218112 694164 220084 694192
rect 218112 694152 218118 694164
rect 220078 694152 220084 694164
rect 220136 694152 220142 694204
rect 457438 694152 457444 694204
rect 457496 694192 457502 694204
rect 462314 694192 462320 694204
rect 457496 694164 462320 694192
rect 457496 694152 457502 694164
rect 462314 694152 462320 694164
rect 462372 694152 462378 694204
rect 504910 694152 504916 694204
rect 504968 694192 504974 694204
rect 510614 694192 510620 694204
rect 504968 694164 510620 694192
rect 504968 694152 504974 694164
rect 510614 694152 510620 694164
rect 510672 694152 510678 694204
rect 552382 694152 552388 694204
rect 552440 694192 552446 694204
rect 558914 694192 558920 694204
rect 552440 694164 558920 694192
rect 552440 694152 552446 694164
rect 558914 694152 558920 694164
rect 558972 694152 558978 694204
rect 578326 672936 578332 672988
rect 578384 672976 578390 672988
rect 580258 672976 580264 672988
rect 578384 672948 580264 672976
rect 578384 672936 578390 672948
rect 580258 672936 580264 672948
rect 580316 672936 580322 672988
rect 578510 659404 578516 659456
rect 578568 659444 578574 659456
rect 580258 659444 580264 659456
rect 578568 659416 580264 659444
rect 578568 659404 578574 659416
rect 580258 659404 580264 659416
rect 580316 659404 580322 659456
rect 578326 646960 578332 647012
rect 578384 647000 578390 647012
rect 580258 647000 580264 647012
rect 578384 646972 580264 647000
rect 578384 646960 578390 646972
rect 580258 646960 580264 646972
rect 580316 646960 580322 647012
rect 578326 620916 578332 620968
rect 578384 620956 578390 620968
rect 580258 620956 580264 620968
rect 578384 620928 580264 620956
rect 578384 620916 578390 620928
rect 580258 620916 580264 620928
rect 580316 620916 580322 620968
rect 578234 510620 578240 510672
rect 578292 510660 578298 510672
rect 580534 510660 580540 510672
rect 578292 510632 580540 510660
rect 578292 510620 578298 510632
rect 580534 510620 580540 510632
rect 580592 510620 580598 510672
rect 578234 470976 578240 471028
rect 578292 471016 578298 471028
rect 579798 471016 579804 471028
rect 578292 470988 579804 471016
rect 578292 470976 578298 470988
rect 579798 470976 579804 470988
rect 579856 470976 579862 471028
rect 578234 404336 578240 404388
rect 578292 404376 578298 404388
rect 580350 404376 580356 404388
rect 578292 404348 580356 404376
rect 578292 404336 578298 404348
rect 580350 404336 580356 404348
rect 580408 404336 580414 404388
rect 578326 362720 578332 362772
rect 578384 362760 578390 362772
rect 580902 362760 580908 362772
rect 578384 362732 580908 362760
rect 578384 362720 578390 362732
rect 580902 362720 580908 362732
rect 580960 362720 580966 362772
rect 578510 219716 578516 219768
rect 578568 219756 578574 219768
rect 580902 219756 580908 219768
rect 578568 219728 580908 219756
rect 578568 219716 578574 219728
rect 580902 219716 580908 219728
rect 580960 219716 580966 219768
rect 578326 181296 578332 181348
rect 578384 181336 578390 181348
rect 580534 181336 580540 181348
rect 578384 181308 580540 181336
rect 578384 181296 578390 181308
rect 580534 181296 580540 181308
rect 580592 181296 580598 181348
rect 578786 142536 578792 142588
rect 578844 142576 578850 142588
rect 580718 142576 580724 142588
rect 578844 142548 580724 142576
rect 578844 142536 578850 142548
rect 580718 142536 580724 142548
rect 580776 142536 580782 142588
rect 578326 116696 578332 116748
rect 578384 116736 578390 116748
rect 580258 116736 580264 116748
rect 578384 116708 580264 116736
rect 578384 116696 578390 116708
rect 580258 116696 580264 116708
rect 580316 116696 580322 116748
rect 578234 60664 578240 60716
rect 578292 60704 578298 60716
rect 580810 60704 580816 60716
rect 578292 60676 580816 60704
rect 578292 60664 578298 60676
rect 580810 60664 580816 60676
rect 580868 60664 580874 60716
rect 578234 20612 578240 20664
rect 578292 20652 578298 20664
rect 580626 20652 580632 20664
rect 578292 20624 580632 20652
rect 578292 20612 578298 20624
rect 580626 20612 580632 20624
rect 580684 20612 580690 20664
rect 1670 4088 1676 4140
rect 1728 4128 1734 4140
rect 20254 4128 20260 4140
rect 1728 4100 20260 4128
rect 1728 4088 1734 4100
rect 20254 4088 20260 4100
rect 20312 4088 20318 4140
rect 21818 4088 21824 4140
rect 21876 4128 21882 4140
rect 39022 4128 39028 4140
rect 21876 4100 39028 4128
rect 21876 4088 21882 4100
rect 39022 4088 39028 4100
rect 39080 4088 39086 4140
rect 43070 4088 43076 4140
rect 43128 4128 43134 4140
rect 58894 4128 58900 4140
rect 43128 4100 58900 4128
rect 43128 4088 43134 4100
rect 58894 4088 58900 4100
rect 58952 4088 58958 4140
rect 66714 4088 66720 4140
rect 66772 4128 66778 4140
rect 80974 4128 80980 4140
rect 66772 4100 80980 4128
rect 66772 4088 66778 4100
rect 80974 4088 80980 4100
rect 81032 4088 81038 4140
rect 83274 4088 83280 4140
rect 83332 4128 83338 4140
rect 96430 4128 96436 4140
rect 83332 4100 96436 4128
rect 83332 4088 83338 4100
rect 96430 4088 96436 4100
rect 96488 4088 96494 4140
rect 97442 4088 97448 4140
rect 97500 4128 97506 4140
rect 109678 4128 109684 4140
rect 97500 4100 109684 4128
rect 97500 4088 97506 4100
rect 109678 4088 109684 4100
rect 109736 4088 109742 4140
rect 112806 4088 112812 4140
rect 112864 4128 112870 4140
rect 124030 4128 124036 4140
rect 112864 4100 124036 4128
rect 112864 4088 112870 4100
rect 124030 4088 124036 4100
rect 124088 4088 124094 4140
rect 124674 4088 124680 4140
rect 124732 4128 124738 4140
rect 135070 4128 135076 4140
rect 124732 4100 135076 4128
rect 124732 4088 124738 4100
rect 135070 4088 135076 4100
rect 135128 4088 135134 4140
rect 136450 4088 136456 4140
rect 136508 4128 136514 4140
rect 146110 4128 146116 4140
rect 136508 4100 146116 4128
rect 136508 4088 136514 4100
rect 146110 4088 146116 4100
rect 146168 4088 146174 4140
rect 157794 4088 157800 4140
rect 157852 4128 157858 4140
rect 165982 4128 165988 4140
rect 157852 4100 165988 4128
rect 157852 4088 157858 4100
rect 165982 4088 165988 4100
rect 166040 4088 166046 4140
rect 174262 4088 174268 4140
rect 174320 4128 174326 4140
rect 181438 4128 181444 4140
rect 174320 4100 181444 4128
rect 174320 4088 174326 4100
rect 181438 4088 181444 4100
rect 181496 4088 181502 4140
rect 415486 4088 415492 4140
rect 415544 4128 415550 4140
rect 424962 4128 424968 4140
rect 415544 4100 424968 4128
rect 415544 4088 415550 4100
rect 424962 4088 424968 4100
rect 425020 4088 425026 4140
rect 430942 4088 430948 4140
rect 431000 4128 431006 4140
rect 441522 4128 441528 4140
rect 431000 4100 441528 4128
rect 431000 4088 431006 4100
rect 441522 4088 441528 4100
rect 441580 4088 441586 4140
rect 464062 4088 464068 4140
rect 464120 4128 464126 4140
rect 476942 4128 476948 4140
rect 464120 4100 476948 4128
rect 464120 4088 464126 4100
rect 476942 4088 476948 4100
rect 477000 4088 477006 4140
rect 477310 4088 477316 4140
rect 477368 4128 477374 4140
rect 491110 4128 491116 4140
rect 477368 4100 491116 4128
rect 477368 4088 477374 4100
rect 491110 4088 491116 4100
rect 491168 4088 491174 4140
rect 493870 4088 493876 4140
rect 493928 4128 493934 4140
rect 508866 4128 508872 4140
rect 493928 4100 508872 4128
rect 493928 4088 493934 4100
rect 508866 4088 508872 4100
rect 508924 4088 508930 4140
rect 510430 4088 510436 4140
rect 510488 4128 510494 4140
rect 525794 4128 525800 4140
rect 510488 4100 525800 4128
rect 510488 4088 510494 4100
rect 525794 4088 525800 4100
rect 525852 4088 525858 4140
rect 525886 4088 525892 4140
rect 525944 4128 525950 4140
rect 543182 4128 543188 4140
rect 525944 4100 543188 4128
rect 525944 4088 525950 4100
rect 543182 4088 543188 4100
rect 543240 4088 543246 4140
rect 549070 4088 549076 4140
rect 549128 4128 549134 4140
rect 568022 4128 568028 4140
rect 549128 4100 568028 4128
rect 549128 4088 549134 4100
rect 568022 4088 568028 4100
rect 568080 4088 568086 4140
rect 15930 4020 15936 4072
rect 15988 4060 15994 4072
rect 33502 4060 33508 4072
rect 15988 4032 33508 4060
rect 15988 4020 15994 4032
rect 33502 4020 33508 4032
rect 33560 4020 33566 4072
rect 40678 4020 40684 4072
rect 40736 4060 40742 4072
rect 56686 4060 56692 4072
rect 40736 4032 56692 4060
rect 40736 4020 40742 4032
rect 56686 4020 56692 4032
rect 56744 4020 56750 4072
rect 62022 4020 62028 4072
rect 62080 4060 62086 4072
rect 76558 4060 76564 4072
rect 62080 4032 76564 4060
rect 62080 4020 62086 4032
rect 76558 4020 76564 4032
rect 76616 4020 76622 4072
rect 77386 4020 77392 4072
rect 77444 4060 77450 4072
rect 90910 4060 90916 4072
rect 77444 4032 90916 4060
rect 77444 4020 77450 4032
rect 90910 4020 90916 4032
rect 90968 4020 90974 4072
rect 93946 4020 93952 4072
rect 94004 4060 94010 4072
rect 106366 4060 106372 4072
rect 94004 4032 106372 4060
rect 94004 4020 94010 4032
rect 106366 4020 106372 4032
rect 106424 4020 106430 4072
rect 119890 4020 119896 4072
rect 119948 4060 119954 4072
rect 130654 4060 130660 4072
rect 119948 4032 130660 4060
rect 119948 4020 119954 4032
rect 130654 4020 130660 4032
rect 130712 4020 130718 4072
rect 132954 4020 132960 4072
rect 133012 4060 133018 4072
rect 142798 4060 142804 4072
rect 133012 4032 142804 4060
rect 133012 4020 133018 4032
rect 142798 4020 142804 4032
rect 142856 4020 142862 4072
rect 143534 4020 143540 4072
rect 143592 4060 143598 4072
rect 152734 4060 152740 4072
rect 143592 4032 152740 4060
rect 143592 4020 143598 4032
rect 152734 4020 152740 4032
rect 152792 4020 152798 4072
rect 154206 4020 154212 4072
rect 154264 4060 154270 4072
rect 162670 4060 162676 4072
rect 154264 4032 162676 4060
rect 154264 4020 154270 4032
rect 162670 4020 162676 4032
rect 162728 4020 162734 4072
rect 168374 4020 168380 4072
rect 168432 4060 168438 4072
rect 175918 4060 175924 4072
rect 168432 4032 175924 4060
rect 168432 4020 168438 4032
rect 175918 4020 175924 4032
rect 175976 4020 175982 4072
rect 176654 4020 176660 4072
rect 176712 4060 176718 4072
rect 183646 4060 183652 4072
rect 176712 4032 183652 4060
rect 176712 4020 176718 4032
rect 183646 4020 183652 4032
rect 183704 4020 183710 4072
rect 400030 4020 400036 4072
rect 400088 4060 400094 4072
rect 408402 4060 408408 4072
rect 400088 4032 408408 4060
rect 400088 4020 400094 4032
rect 408402 4020 408408 4032
rect 408460 4020 408466 4072
rect 421006 4020 421012 4072
rect 421064 4060 421070 4072
rect 430850 4060 430856 4072
rect 421064 4032 430856 4060
rect 421064 4020 421070 4032
rect 430850 4020 430856 4032
rect 430908 4020 430914 4072
rect 432046 4020 432052 4072
rect 432104 4060 432110 4072
rect 442626 4060 442632 4072
rect 432104 4032 442632 4060
rect 432104 4020 432110 4032
rect 442626 4020 442632 4032
rect 442684 4020 442690 4072
rect 448606 4020 448612 4072
rect 448664 4060 448670 4072
rect 460382 4060 460388 4072
rect 448664 4032 460388 4060
rect 448664 4020 448670 4032
rect 460382 4020 460388 4032
rect 460440 4020 460446 4072
rect 465166 4020 465172 4072
rect 465224 4060 465230 4072
rect 465224 4032 476160 4060
rect 465224 4020 465230 4032
rect 6454 3952 6460 4004
rect 6512 3992 6518 4004
rect 24670 3992 24676 4004
rect 6512 3964 24676 3992
rect 6512 3952 6518 3964
rect 24670 3952 24676 3964
rect 24728 3952 24734 4004
rect 39574 3952 39580 4004
rect 39632 3992 39638 4004
rect 55582 3992 55588 4004
rect 39632 3964 55588 3992
rect 39632 3952 39638 3964
rect 55582 3952 55588 3964
rect 55640 3952 55646 4004
rect 58434 3952 58440 4004
rect 58492 3992 58498 4004
rect 73246 3992 73252 4004
rect 58492 3964 73252 3992
rect 58492 3952 58498 3964
rect 73246 3952 73252 3964
rect 73304 3952 73310 4004
rect 84470 3952 84476 4004
rect 84528 3992 84534 4004
rect 97534 3992 97540 4004
rect 84528 3964 97540 3992
rect 84528 3952 84534 3964
rect 97534 3952 97540 3964
rect 97592 3952 97598 4004
rect 101030 3952 101036 4004
rect 101088 3992 101094 4004
rect 112990 3992 112996 4004
rect 101088 3964 112996 3992
rect 101088 3952 101094 3964
rect 112990 3952 112996 3964
rect 113048 3952 113054 4004
rect 115290 3952 115296 4004
rect 115348 3992 115354 4004
rect 126238 3992 126244 4004
rect 115348 3964 126244 3992
rect 115348 3952 115354 3964
rect 126238 3952 126244 3964
rect 126296 3952 126302 4004
rect 126974 3952 126980 4004
rect 127032 3992 127038 4004
rect 137278 3992 137284 4004
rect 127032 3964 137284 3992
rect 127032 3952 127038 3964
rect 137278 3952 137284 3964
rect 137336 3952 137342 4004
rect 150618 3952 150624 4004
rect 150676 3992 150682 4004
rect 159358 3992 159364 4004
rect 150676 3964 159364 3992
rect 150676 3952 150682 3964
rect 159358 3952 159364 3964
rect 159416 3952 159422 4004
rect 180242 3952 180248 4004
rect 180300 3992 180306 4004
rect 186958 3992 186964 4004
rect 180300 3964 186964 3992
rect 180300 3952 180306 3964
rect 186958 3952 186964 3964
rect 187016 3952 187022 4004
rect 189718 3952 189724 4004
rect 189776 3992 189782 4004
rect 195790 3992 195796 4004
rect 189776 3964 195796 3992
rect 189776 3952 189782 3964
rect 195790 3952 195796 3964
rect 195848 3952 195854 4004
rect 407758 3952 407764 4004
rect 407816 3992 407822 4004
rect 407816 3964 416544 3992
rect 407816 3952 407822 3964
rect 13538 3884 13544 3936
rect 13596 3924 13602 3936
rect 31294 3924 31300 3936
rect 13596 3896 31300 3924
rect 13596 3884 13602 3896
rect 31294 3884 31300 3896
rect 31352 3884 31358 3936
rect 38378 3884 38384 3936
rect 38436 3924 38442 3936
rect 54478 3924 54484 3936
rect 38436 3896 54484 3924
rect 38436 3884 38442 3896
rect 54478 3884 54484 3896
rect 54536 3884 54542 3936
rect 57238 3884 57244 3936
rect 57296 3924 57302 3936
rect 72142 3924 72148 3936
rect 57296 3896 72148 3924
rect 57296 3884 57302 3896
rect 72142 3884 72148 3896
rect 72200 3884 72206 3936
rect 78582 3884 78588 3936
rect 78640 3924 78646 3936
rect 92014 3924 92020 3936
rect 78640 3896 92020 3924
rect 78640 3884 78646 3896
rect 92014 3884 92020 3896
rect 92072 3884 92078 3936
rect 92750 3884 92756 3936
rect 92808 3924 92814 3936
rect 105262 3924 105268 3936
rect 92808 3896 105268 3924
rect 92808 3884 92814 3896
rect 105262 3884 105268 3896
rect 105320 3884 105326 3936
rect 108114 3884 108120 3936
rect 108172 3924 108178 3936
rect 119614 3924 119620 3936
rect 108172 3896 119620 3924
rect 108172 3884 108178 3896
rect 119614 3884 119620 3896
rect 119672 3884 119678 3936
rect 122282 3884 122288 3936
rect 122340 3924 122346 3936
rect 132862 3924 132868 3936
rect 122340 3896 132868 3924
rect 122340 3884 122346 3896
rect 132862 3884 132868 3896
rect 132920 3884 132926 3936
rect 134150 3884 134156 3936
rect 134208 3924 134214 3936
rect 143902 3924 143908 3936
rect 134208 3896 143908 3924
rect 134208 3884 134214 3896
rect 143902 3884 143908 3896
rect 143960 3884 143966 3936
rect 149514 3884 149520 3936
rect 149572 3924 149578 3936
rect 158254 3924 158260 3936
rect 149572 3896 158260 3924
rect 149572 3884 149578 3896
rect 158254 3884 158260 3896
rect 158312 3884 158318 3936
rect 160094 3884 160100 3936
rect 160152 3924 160158 3936
rect 168190 3924 168196 3936
rect 160152 3896 168196 3924
rect 160152 3884 160158 3896
rect 168190 3884 168196 3896
rect 168248 3884 168254 3936
rect 179046 3884 179052 3936
rect 179104 3924 179110 3936
rect 185854 3924 185860 3936
rect 179104 3896 185860 3924
rect 179104 3884 179110 3896
rect 185854 3884 185860 3896
rect 185912 3884 185918 3936
rect 401134 3884 401140 3936
rect 401192 3924 401198 3936
rect 401192 3896 408816 3924
rect 401192 3884 401198 3896
rect 8754 3816 8760 3868
rect 8812 3856 8818 3868
rect 26878 3856 26884 3868
rect 8812 3828 26884 3856
rect 8812 3816 8818 3828
rect 26878 3816 26884 3828
rect 26936 3816 26942 3868
rect 32490 3816 32496 3868
rect 32548 3856 32554 3868
rect 48958 3856 48964 3868
rect 32548 3828 48964 3856
rect 32548 3816 32554 3828
rect 48958 3816 48964 3828
rect 49016 3816 49022 3868
rect 53742 3816 53748 3868
rect 53800 3856 53806 3868
rect 68830 3856 68836 3868
rect 53800 3828 68836 3856
rect 53800 3816 53806 3828
rect 68830 3816 68836 3828
rect 68888 3816 68894 3868
rect 71498 3816 71504 3868
rect 71556 3856 71562 3868
rect 85390 3856 85396 3868
rect 71556 3828 85396 3856
rect 71556 3816 71562 3828
rect 85390 3816 85396 3828
rect 85448 3816 85454 3868
rect 89162 3816 89168 3868
rect 89220 3856 89226 3868
rect 101950 3856 101956 3868
rect 89220 3828 101956 3856
rect 89220 3816 89226 3828
rect 101950 3816 101956 3828
rect 102008 3816 102014 3868
rect 103330 3816 103336 3868
rect 103388 3856 103394 3868
rect 115198 3856 115204 3868
rect 103388 3828 115204 3856
rect 103388 3816 103394 3828
rect 115198 3816 115204 3828
rect 115256 3816 115262 3868
rect 116394 3816 116400 3868
rect 116452 3856 116458 3868
rect 127342 3856 127348 3868
rect 116452 3828 127348 3856
rect 116452 3816 116458 3828
rect 127342 3816 127348 3828
rect 127400 3816 127406 3868
rect 137646 3816 137652 3868
rect 137704 3856 137710 3868
rect 147214 3856 147220 3868
rect 137704 3828 147220 3856
rect 137704 3816 137710 3828
rect 147214 3816 147220 3828
rect 147272 3816 147278 3868
rect 148318 3816 148324 3868
rect 148376 3856 148382 3868
rect 157150 3856 157156 3868
rect 148376 3828 157156 3856
rect 148376 3816 148382 3828
rect 157150 3816 157156 3828
rect 157208 3816 157214 3868
rect 161290 3816 161296 3868
rect 161348 3856 161354 3868
rect 169294 3856 169300 3868
rect 161348 3828 169300 3856
rect 161348 3816 161354 3828
rect 169294 3816 169300 3828
rect 169352 3816 169358 3868
rect 353662 3816 353668 3868
rect 353720 3856 353726 3868
rect 358722 3856 358728 3868
rect 353720 3828 358728 3856
rect 353720 3816 353726 3828
rect 358722 3816 358728 3828
rect 358780 3816 358786 3868
rect 371326 3816 371332 3868
rect 371384 3856 371390 3868
rect 377674 3856 377680 3868
rect 371384 3828 377680 3856
rect 371384 3816 371390 3828
rect 377674 3816 377680 3828
rect 377732 3816 377738 3868
rect 397822 3816 397828 3868
rect 397880 3856 397886 3868
rect 406010 3856 406016 3868
rect 397880 3828 406016 3856
rect 397880 3816 397886 3828
rect 406010 3816 406016 3828
rect 406068 3816 406074 3868
rect 408788 3856 408816 3896
rect 408862 3884 408868 3936
rect 408920 3924 408926 3936
rect 416516 3924 416544 3964
rect 416590 3952 416596 4004
rect 416648 3992 416654 4004
rect 426158 3992 426164 4004
rect 416648 3964 426164 3992
rect 416648 3952 416654 3964
rect 426158 3952 426164 3964
rect 426216 3952 426222 4004
rect 426526 3952 426532 4004
rect 426584 3992 426590 4004
rect 436738 3992 436744 4004
rect 426584 3964 436744 3992
rect 426584 3952 426590 3964
rect 436738 3952 436744 3964
rect 436796 3952 436802 4004
rect 437566 3952 437572 4004
rect 437624 3992 437630 4004
rect 448514 3992 448520 4004
rect 437624 3964 448520 3992
rect 437624 3952 437630 3964
rect 448514 3952 448520 3964
rect 448572 3952 448578 4004
rect 461854 3952 461860 4004
rect 461912 3992 461918 4004
rect 474550 3992 474556 4004
rect 461912 3964 474556 3992
rect 461912 3952 461918 3964
rect 474550 3952 474556 3964
rect 474608 3952 474614 4004
rect 476132 3992 476160 4032
rect 476206 4020 476212 4072
rect 476264 4060 476270 4072
rect 481634 4060 481640 4072
rect 476264 4032 481640 4060
rect 476264 4020 476270 4032
rect 481634 4020 481640 4032
rect 481692 4020 481698 4072
rect 481726 4020 481732 4072
rect 481784 4060 481790 4072
rect 495894 4060 495900 4072
rect 481784 4032 495900 4060
rect 481784 4020 481790 4032
rect 495894 4020 495900 4032
rect 495952 4020 495958 4072
rect 498286 4020 498292 4072
rect 498344 4060 498350 4072
rect 513558 4060 513564 4072
rect 498344 4032 513564 4060
rect 498344 4020 498350 4032
rect 513558 4020 513564 4032
rect 513616 4020 513622 4072
rect 520366 4020 520372 4072
rect 520424 4060 520430 4072
rect 536834 4060 536840 4072
rect 520424 4032 536840 4060
rect 520424 4020 520430 4032
rect 536834 4020 536840 4032
rect 536892 4020 536898 4072
rect 536926 4020 536932 4072
rect 536984 4060 536990 4072
rect 554958 4060 554964 4072
rect 536984 4032 554964 4060
rect 536984 4020 536990 4032
rect 554958 4020 554964 4032
rect 555016 4020 555022 4072
rect 556798 4020 556804 4072
rect 556856 4060 556862 4072
rect 576302 4060 576308 4072
rect 556856 4032 576308 4060
rect 556856 4020 556862 4032
rect 576302 4020 576308 4032
rect 576360 4020 576366 4072
rect 478138 3992 478144 4004
rect 476132 3964 478144 3992
rect 478138 3952 478144 3964
rect 478196 3952 478202 4004
rect 478414 3952 478420 4004
rect 478472 3992 478478 4004
rect 492306 3992 492312 4004
rect 478472 3964 492312 3992
rect 478472 3952 478478 3964
rect 492306 3952 492312 3964
rect 492364 3952 492370 4004
rect 497182 3952 497188 4004
rect 497240 3992 497246 4004
rect 512454 3992 512460 4004
rect 497240 3964 512460 3992
rect 497240 3952 497246 3964
rect 512454 3952 512460 3964
rect 512512 3952 512518 4004
rect 513742 3952 513748 4004
rect 513800 3992 513806 4004
rect 530118 3992 530124 4004
rect 513800 3964 530124 3992
rect 513800 3952 513806 3964
rect 530118 3952 530124 3964
rect 530176 3952 530182 4004
rect 530302 3952 530308 4004
rect 530360 3992 530366 4004
rect 547874 3992 547880 4004
rect 530360 3964 547880 3992
rect 530360 3952 530366 3964
rect 547874 3952 547880 3964
rect 547932 3952 547938 4004
rect 550174 3952 550180 4004
rect 550232 3992 550238 4004
rect 569126 3992 569132 4004
rect 550232 3964 569132 3992
rect 550232 3952 550238 3964
rect 569126 3952 569132 3964
rect 569184 3952 569190 4004
rect 416682 3924 416688 3936
rect 408920 3896 416360 3924
rect 416516 3896 416688 3924
rect 408920 3884 408926 3896
rect 409598 3856 409604 3868
rect 408788 3828 409604 3856
rect 409598 3816 409604 3828
rect 409656 3816 409662 3868
rect 409966 3816 409972 3868
rect 410024 3856 410030 3868
rect 416332 3856 416360 3896
rect 416682 3884 416688 3896
rect 416740 3884 416746 3936
rect 417694 3884 417700 3936
rect 417752 3924 417758 3936
rect 427262 3924 427268 3936
rect 417752 3896 427268 3924
rect 417752 3884 417758 3896
rect 427262 3884 427268 3896
rect 427320 3884 427326 3936
rect 427630 3884 427636 3936
rect 427688 3924 427694 3936
rect 437934 3924 437940 3936
rect 427688 3896 437940 3924
rect 427688 3884 427694 3896
rect 437934 3884 437940 3896
rect 437992 3884 437998 3936
rect 441982 3884 441988 3936
rect 442040 3924 442046 3936
rect 453298 3924 453304 3936
rect 442040 3896 453304 3924
rect 442040 3884 442046 3896
rect 453298 3884 453304 3896
rect 453356 3884 453362 3936
rect 457438 3884 457444 3936
rect 457496 3924 457502 3936
rect 469858 3924 469864 3936
rect 457496 3896 469864 3924
rect 457496 3884 457502 3896
rect 469858 3884 469864 3896
rect 469916 3884 469922 3936
rect 471790 3884 471796 3936
rect 471848 3924 471854 3936
rect 485222 3924 485228 3936
rect 471848 3896 485228 3924
rect 471848 3884 471854 3896
rect 485222 3884 485228 3896
rect 485280 3884 485286 3936
rect 488350 3884 488356 3936
rect 488408 3924 488414 3936
rect 488408 3896 502656 3924
rect 488408 3884 488414 3896
rect 417878 3856 417884 3868
rect 410024 3828 416268 3856
rect 416332 3828 417884 3856
rect 410024 3816 410030 3828
rect 566 3748 572 3800
rect 624 3788 630 3800
rect 19150 3788 19156 3800
rect 624 3760 19156 3788
rect 624 3748 630 3760
rect 19150 3748 19156 3760
rect 19208 3748 19214 3800
rect 23014 3748 23020 3800
rect 23072 3788 23078 3800
rect 40126 3788 40132 3800
rect 23072 3760 40132 3788
rect 23072 3748 23078 3760
rect 40126 3748 40132 3760
rect 40184 3748 40190 3800
rect 41874 3748 41880 3800
rect 41932 3788 41938 3800
rect 57790 3788 57796 3800
rect 41932 3760 57796 3788
rect 41932 3748 41938 3760
rect 57790 3748 57796 3760
rect 57848 3748 57854 3800
rect 63218 3748 63224 3800
rect 63276 3788 63282 3800
rect 77662 3788 77668 3800
rect 63276 3760 77668 3788
rect 63276 3748 63282 3760
rect 77662 3748 77668 3760
rect 77720 3748 77726 3800
rect 79686 3748 79692 3800
rect 79744 3788 79750 3800
rect 93118 3788 93124 3800
rect 79744 3760 93124 3788
rect 79744 3748 79750 3760
rect 93118 3748 93124 3760
rect 93176 3748 93182 3800
rect 96246 3748 96252 3800
rect 96304 3788 96310 3800
rect 108574 3788 108580 3800
rect 96304 3760 108580 3788
rect 96304 3748 96310 3760
rect 108574 3748 108580 3760
rect 108632 3748 108638 3800
rect 110506 3748 110512 3800
rect 110564 3788 110570 3800
rect 121822 3788 121828 3800
rect 110564 3760 121828 3788
rect 110564 3748 110570 3760
rect 121822 3748 121828 3760
rect 121880 3748 121886 3800
rect 123478 3748 123484 3800
rect 123536 3788 123542 3800
rect 133966 3788 133972 3800
rect 123536 3760 133972 3788
rect 123536 3748 123542 3760
rect 133966 3748 133972 3760
rect 134024 3748 134030 3800
rect 140038 3748 140044 3800
rect 140096 3788 140102 3800
rect 149422 3788 149428 3800
rect 140096 3760 149428 3788
rect 140096 3748 140102 3760
rect 149422 3748 149428 3760
rect 149480 3748 149486 3800
rect 167178 3748 167184 3800
rect 167236 3788 167242 3800
rect 174814 3788 174820 3800
rect 167236 3760 174820 3788
rect 167236 3748 167242 3760
rect 174814 3748 174820 3760
rect 174872 3748 174878 3800
rect 175458 3748 175464 3800
rect 175516 3788 175522 3800
rect 182542 3788 182548 3800
rect 175516 3760 182548 3788
rect 175516 3748 175522 3760
rect 182542 3748 182548 3760
rect 182600 3748 182606 3800
rect 197906 3748 197912 3800
rect 197964 3788 197970 3800
rect 203518 3788 203524 3800
rect 197964 3760 203524 3788
rect 197964 3748 197970 3760
rect 203518 3748 203524 3760
rect 203576 3748 203582 3800
rect 208578 3748 208584 3800
rect 208636 3788 208642 3800
rect 213454 3788 213460 3800
rect 208636 3760 213460 3788
rect 208636 3748 208642 3760
rect 213454 3748 213460 3760
rect 213512 3748 213518 3800
rect 218054 3748 218060 3800
rect 218112 3788 218118 3800
rect 222286 3788 222292 3800
rect 218112 3760 222292 3788
rect 218112 3748 218118 3760
rect 222286 3748 222292 3760
rect 222344 3748 222350 3800
rect 381262 3748 381268 3800
rect 381320 3788 381326 3800
rect 388254 3788 388260 3800
rect 381320 3760 388260 3788
rect 381320 3748 381326 3760
rect 388254 3748 388260 3760
rect 388312 3748 388318 3800
rect 398926 3748 398932 3800
rect 398984 3788 398990 3800
rect 407206 3788 407212 3800
rect 398984 3760 407212 3788
rect 398984 3748 398990 3760
rect 407206 3748 407212 3760
rect 407264 3748 407270 3800
rect 411070 3748 411076 3800
rect 411128 3788 411134 3800
rect 416240 3788 416268 3828
rect 417878 3816 417884 3828
rect 417936 3816 417942 3868
rect 424318 3816 424324 3868
rect 424376 3856 424382 3868
rect 434438 3856 434444 3868
rect 424376 3828 434444 3856
rect 424376 3816 424382 3828
rect 434438 3816 434444 3828
rect 434496 3816 434502 3868
rect 434530 3816 434536 3868
rect 434588 3856 434594 3868
rect 445018 3856 445024 3868
rect 434588 3828 445024 3856
rect 434588 3816 434594 3828
rect 445018 3816 445024 3828
rect 445076 3816 445082 3868
rect 446398 3816 446404 3868
rect 446456 3856 446462 3868
rect 458082 3856 458088 3868
rect 446456 3828 458088 3856
rect 446456 3816 446462 3828
rect 458082 3816 458088 3828
rect 458140 3816 458146 3868
rect 458542 3816 458548 3868
rect 458600 3856 458606 3868
rect 471054 3856 471060 3868
rect 458600 3828 471060 3856
rect 458600 3816 458606 3828
rect 471054 3816 471060 3828
rect 471112 3816 471118 3868
rect 473998 3816 474004 3868
rect 474056 3856 474062 3868
rect 487614 3856 487620 3868
rect 474056 3828 487620 3856
rect 474056 3816 474062 3828
rect 487614 3816 487620 3828
rect 487672 3816 487678 3868
rect 497090 3856 497096 3868
rect 489886 3828 497096 3856
rect 418982 3788 418988 3800
rect 411128 3760 412634 3788
rect 416240 3760 418988 3788
rect 411128 3748 411134 3760
rect 9950 3680 9956 3732
rect 10008 3720 10014 3732
rect 27982 3720 27988 3732
rect 10008 3692 27988 3720
rect 10008 3680 10014 3692
rect 27982 3680 27988 3692
rect 28040 3680 28046 3732
rect 31294 3680 31300 3732
rect 31352 3720 31358 3732
rect 47854 3720 47860 3732
rect 31352 3692 47860 3720
rect 31352 3680 31358 3692
rect 47854 3680 47860 3692
rect 47912 3680 47918 3732
rect 50154 3680 50160 3732
rect 50212 3720 50218 3732
rect 65518 3720 65524 3732
rect 50212 3692 65524 3720
rect 50212 3680 50218 3692
rect 65518 3680 65524 3692
rect 65576 3680 65582 3732
rect 74994 3680 75000 3732
rect 75052 3720 75058 3732
rect 88702 3720 88708 3732
rect 75052 3692 88708 3720
rect 75052 3680 75058 3692
rect 88702 3680 88708 3692
rect 88760 3680 88766 3732
rect 91554 3680 91560 3732
rect 91612 3720 91618 3732
rect 104158 3720 104164 3732
rect 91612 3692 104164 3720
rect 91612 3680 91618 3692
rect 104158 3680 104164 3692
rect 104216 3680 104222 3732
rect 117590 3680 117596 3732
rect 117648 3720 117654 3732
rect 128446 3720 128452 3732
rect 117648 3692 128452 3720
rect 117648 3680 117654 3692
rect 128446 3680 128452 3692
rect 128504 3680 128510 3732
rect 138842 3680 138848 3732
rect 138900 3720 138906 3732
rect 147950 3720 147956 3732
rect 138900 3692 147956 3720
rect 138900 3680 138906 3692
rect 147950 3680 147956 3692
rect 148008 3680 148014 3732
rect 177850 3680 177856 3732
rect 177908 3720 177914 3732
rect 184750 3720 184756 3732
rect 177908 3692 184756 3720
rect 177908 3680 177914 3692
rect 184750 3680 184756 3692
rect 184808 3680 184814 3732
rect 228726 3680 228732 3732
rect 228784 3720 228790 3732
rect 232222 3720 232228 3732
rect 228784 3692 232228 3720
rect 228784 3680 228790 3692
rect 232222 3680 232228 3692
rect 232280 3680 232286 3732
rect 412606 3720 412634 3760
rect 418982 3748 418988 3760
rect 419040 3748 419046 3800
rect 423214 3748 423220 3800
rect 423272 3788 423278 3800
rect 433242 3788 433248 3800
rect 423272 3760 433248 3788
rect 423272 3748 423278 3760
rect 433242 3748 433248 3760
rect 433300 3748 433306 3800
rect 435358 3748 435364 3800
rect 435416 3788 435422 3800
rect 446214 3788 446220 3800
rect 435416 3760 446220 3788
rect 435416 3748 435422 3760
rect 446214 3748 446220 3760
rect 446272 3748 446278 3800
rect 451918 3748 451924 3800
rect 451976 3788 451982 3800
rect 463970 3788 463976 3800
rect 451976 3760 463976 3788
rect 451976 3748 451982 3760
rect 463970 3748 463976 3760
rect 464028 3748 464034 3800
rect 467374 3748 467380 3800
rect 467432 3788 467438 3800
rect 475378 3788 475384 3800
rect 467432 3760 475384 3788
rect 467432 3748 467438 3760
rect 475378 3748 475384 3760
rect 475436 3748 475442 3800
rect 482830 3748 482836 3800
rect 482888 3788 482894 3800
rect 489886 3788 489914 3828
rect 497090 3816 497096 3828
rect 497148 3816 497154 3868
rect 502628 3856 502656 3896
rect 502702 3884 502708 3936
rect 502760 3924 502766 3936
rect 517974 3924 517980 3936
rect 502760 3896 517980 3924
rect 502760 3884 502766 3896
rect 517974 3884 517980 3896
rect 518032 3884 518038 3936
rect 518158 3884 518164 3936
rect 518216 3924 518222 3936
rect 534534 3924 534540 3936
rect 518216 3896 534540 3924
rect 518216 3884 518222 3896
rect 534534 3884 534540 3896
rect 534592 3884 534598 3936
rect 534718 3884 534724 3936
rect 534776 3924 534782 3936
rect 552658 3924 552664 3936
rect 534776 3896 552664 3924
rect 534776 3884 534782 3896
rect 552658 3884 552664 3896
rect 552716 3884 552722 3936
rect 553486 3884 553492 3936
rect 553544 3924 553550 3936
rect 572714 3924 572720 3936
rect 553544 3896 572720 3924
rect 553544 3884 553550 3896
rect 572714 3884 572720 3896
rect 572772 3884 572778 3936
rect 502978 3856 502984 3868
rect 502628 3828 502984 3856
rect 502978 3816 502984 3828
rect 503036 3816 503042 3868
rect 506474 3856 506480 3868
rect 504836 3828 506480 3856
rect 482888 3760 489914 3788
rect 482888 3748 482894 3760
rect 491662 3748 491668 3800
rect 491720 3788 491726 3800
rect 504836 3788 504864 3828
rect 506474 3816 506480 3828
rect 506532 3816 506538 3868
rect 514846 3816 514852 3868
rect 514904 3856 514910 3868
rect 531314 3856 531320 3868
rect 514904 3828 531320 3856
rect 514904 3816 514910 3828
rect 531314 3816 531320 3828
rect 531372 3816 531378 3868
rect 533614 3816 533620 3868
rect 533672 3856 533678 3868
rect 551094 3856 551100 3868
rect 533672 3828 551100 3856
rect 533672 3816 533678 3828
rect 551094 3816 551100 3828
rect 551152 3816 551158 3868
rect 551278 3816 551284 3868
rect 551336 3856 551342 3868
rect 570322 3856 570328 3868
rect 551336 3828 570328 3856
rect 551336 3816 551342 3828
rect 570322 3816 570328 3828
rect 570380 3816 570386 3868
rect 491720 3760 504864 3788
rect 491720 3748 491726 3760
rect 504910 3748 504916 3800
rect 504968 3788 504974 3800
rect 520734 3788 520740 3800
rect 504968 3760 520740 3788
rect 504968 3748 504974 3760
rect 520734 3748 520740 3760
rect 520792 3748 520798 3800
rect 529198 3748 529204 3800
rect 529256 3788 529262 3800
rect 546678 3788 546684 3800
rect 529256 3760 546684 3788
rect 529256 3748 529262 3760
rect 546678 3748 546684 3760
rect 546736 3748 546742 3800
rect 557902 3748 557908 3800
rect 557960 3788 557966 3800
rect 577406 3788 577412 3800
rect 557960 3760 577412 3788
rect 557960 3748 557966 3760
rect 577406 3748 577412 3760
rect 577464 3748 577470 3800
rect 420178 3720 420184 3732
rect 412606 3692 420184 3720
rect 420178 3680 420184 3692
rect 420236 3680 420242 3732
rect 423766 3720 423772 3732
rect 420288 3692 423772 3720
rect 14734 3612 14740 3664
rect 14792 3652 14798 3664
rect 32398 3652 32404 3664
rect 14792 3624 32404 3652
rect 14792 3612 14798 3624
rect 32398 3612 32404 3624
rect 32456 3612 32462 3664
rect 34790 3612 34796 3664
rect 34848 3652 34854 3664
rect 51166 3652 51172 3664
rect 34848 3624 51172 3652
rect 34848 3612 34854 3624
rect 51166 3612 51172 3624
rect 51224 3612 51230 3664
rect 56042 3612 56048 3664
rect 56100 3652 56106 3664
rect 71038 3652 71044 3664
rect 56100 3624 71044 3652
rect 56100 3612 56106 3624
rect 71038 3612 71044 3624
rect 71096 3612 71102 3664
rect 82078 3612 82084 3664
rect 82136 3652 82142 3664
rect 95326 3652 95332 3664
rect 82136 3624 95332 3652
rect 82136 3612 82142 3624
rect 95326 3612 95332 3624
rect 95384 3612 95390 3664
rect 99834 3612 99840 3664
rect 99892 3652 99898 3664
rect 111886 3652 111892 3664
rect 99892 3624 111892 3652
rect 99892 3612 99898 3624
rect 111886 3612 111892 3624
rect 111944 3612 111950 3664
rect 114002 3612 114008 3664
rect 114060 3652 114066 3664
rect 125134 3652 125140 3664
rect 114060 3624 125140 3652
rect 114060 3612 114066 3624
rect 125134 3612 125140 3624
rect 125192 3612 125198 3664
rect 131758 3612 131764 3664
rect 131816 3652 131822 3664
rect 141694 3652 141700 3664
rect 131816 3624 141700 3652
rect 131816 3612 131822 3624
rect 141694 3612 141700 3624
rect 141752 3612 141758 3664
rect 144730 3612 144736 3664
rect 144788 3652 144794 3664
rect 153838 3652 153844 3664
rect 144788 3624 153844 3652
rect 144788 3612 144794 3624
rect 153838 3612 153844 3624
rect 153896 3612 153902 3664
rect 343726 3612 343732 3664
rect 343784 3652 343790 3664
rect 348050 3652 348056 3664
rect 343784 3624 348056 3652
rect 343784 3612 343790 3624
rect 348050 3612 348056 3624
rect 348108 3612 348114 3664
rect 363598 3612 363604 3664
rect 363656 3652 363662 3664
rect 369394 3652 369400 3664
rect 363656 3624 369400 3652
rect 363656 3612 363662 3624
rect 369394 3612 369400 3624
rect 369452 3612 369458 3664
rect 380158 3612 380164 3664
rect 380216 3652 380222 3664
rect 387150 3652 387156 3664
rect 380216 3624 387156 3652
rect 380216 3612 380222 3624
rect 387150 3612 387156 3624
rect 387208 3612 387214 3664
rect 391198 3612 391204 3664
rect 391256 3652 391262 3664
rect 398926 3652 398932 3664
rect 391256 3624 398932 3652
rect 391256 3612 391262 3624
rect 398926 3612 398932 3624
rect 398984 3612 398990 3664
rect 405550 3612 405556 3664
rect 405608 3652 405614 3664
rect 414290 3652 414296 3664
rect 405608 3624 414296 3652
rect 405608 3612 405614 3624
rect 414290 3612 414296 3624
rect 414348 3612 414354 3664
rect 414382 3612 414388 3664
rect 414440 3652 414446 3664
rect 420288 3652 420316 3692
rect 423766 3680 423772 3692
rect 423824 3680 423830 3732
rect 425422 3680 425428 3732
rect 425480 3720 425486 3732
rect 435542 3720 435548 3732
rect 425480 3692 435548 3720
rect 425480 3680 425486 3692
rect 435542 3680 435548 3692
rect 435600 3680 435606 3732
rect 436462 3680 436468 3732
rect 436520 3720 436526 3732
rect 447410 3720 447416 3732
rect 436520 3692 447416 3720
rect 436520 3680 436526 3692
rect 447410 3680 447416 3692
rect 447468 3680 447474 3732
rect 450814 3680 450820 3732
rect 450872 3720 450878 3732
rect 462774 3720 462780 3732
rect 450872 3692 462780 3720
rect 450872 3680 450878 3692
rect 462774 3680 462780 3692
rect 462832 3680 462838 3732
rect 462958 3680 462964 3732
rect 463016 3720 463022 3732
rect 474734 3720 474740 3732
rect 463016 3692 474740 3720
rect 463016 3680 463022 3692
rect 474734 3680 474740 3692
rect 474792 3680 474798 3732
rect 475470 3680 475476 3732
rect 475528 3720 475534 3732
rect 488810 3720 488816 3732
rect 475528 3692 488816 3720
rect 475528 3680 475534 3692
rect 488810 3680 488816 3692
rect 488868 3680 488874 3732
rect 494974 3680 494980 3732
rect 495032 3720 495038 3732
rect 510062 3720 510068 3732
rect 495032 3692 510068 3720
rect 495032 3680 495038 3692
rect 510062 3680 510068 3692
rect 510120 3680 510126 3732
rect 511534 3680 511540 3732
rect 511592 3720 511598 3732
rect 527818 3720 527824 3732
rect 511592 3692 527824 3720
rect 511592 3680 511598 3692
rect 527818 3680 527824 3692
rect 527876 3680 527882 3732
rect 528094 3680 528100 3732
rect 528152 3720 528158 3732
rect 545482 3720 545488 3732
rect 528152 3692 545488 3720
rect 528152 3680 528158 3692
rect 545482 3680 545488 3692
rect 545540 3680 545546 3732
rect 545758 3680 545764 3732
rect 545816 3720 545822 3732
rect 564434 3720 564440 3732
rect 545816 3692 564440 3720
rect 545816 3680 545822 3692
rect 564434 3680 564440 3692
rect 564492 3680 564498 3732
rect 429654 3652 429660 3664
rect 414440 3624 420316 3652
rect 421852 3624 429660 3652
rect 414440 3612 414446 3624
rect 11146 3544 11152 3596
rect 11204 3584 11210 3596
rect 29086 3584 29092 3596
rect 11204 3556 29092 3584
rect 11204 3544 11210 3556
rect 29086 3544 29092 3556
rect 29144 3544 29150 3596
rect 46658 3544 46664 3596
rect 46716 3584 46722 3596
rect 62206 3584 62212 3596
rect 46716 3556 62212 3584
rect 46716 3544 46722 3556
rect 62206 3544 62212 3556
rect 62264 3544 62270 3596
rect 64322 3544 64328 3596
rect 64380 3584 64386 3596
rect 78766 3584 78772 3596
rect 64380 3556 78772 3584
rect 64380 3544 64386 3556
rect 78766 3544 78772 3556
rect 78824 3544 78830 3596
rect 80882 3544 80888 3596
rect 80940 3584 80946 3596
rect 94222 3584 94228 3596
rect 80940 3556 94228 3584
rect 80940 3544 80946 3556
rect 94222 3544 94228 3556
rect 94280 3544 94286 3596
rect 98638 3544 98644 3596
rect 98696 3584 98702 3596
rect 110782 3584 110788 3596
rect 98696 3556 110788 3584
rect 98696 3544 98702 3556
rect 110782 3544 110788 3556
rect 110840 3544 110846 3596
rect 111610 3544 111616 3596
rect 111668 3584 111674 3596
rect 122926 3584 122932 3596
rect 111668 3556 122932 3584
rect 111668 3544 111674 3556
rect 122926 3544 122932 3556
rect 122984 3544 122990 3596
rect 128170 3544 128176 3596
rect 128228 3584 128234 3596
rect 138382 3584 138388 3596
rect 128228 3556 138388 3584
rect 128228 3544 128234 3556
rect 138382 3544 138388 3556
rect 138440 3544 138446 3596
rect 145926 3544 145932 3596
rect 145984 3584 145990 3596
rect 154942 3584 154948 3596
rect 145984 3556 154948 3584
rect 145984 3544 145990 3556
rect 154942 3544 154948 3556
rect 155000 3544 155006 3596
rect 156598 3544 156604 3596
rect 156656 3584 156662 3596
rect 164878 3584 164884 3596
rect 156656 3556 164884 3584
rect 156656 3544 156662 3556
rect 164878 3544 164884 3556
rect 164936 3544 164942 3596
rect 169570 3544 169576 3596
rect 169628 3584 169634 3596
rect 177022 3584 177028 3596
rect 169628 3556 177028 3584
rect 169628 3544 169634 3556
rect 177022 3544 177028 3556
rect 177080 3544 177086 3596
rect 193214 3544 193220 3596
rect 193272 3584 193278 3596
rect 199102 3584 199108 3596
rect 193272 3556 199108 3584
rect 193272 3544 193278 3556
rect 199102 3544 199108 3556
rect 199160 3544 199166 3596
rect 334894 3544 334900 3596
rect 334952 3584 334958 3596
rect 338666 3584 338672 3596
rect 334952 3556 338672 3584
rect 334952 3544 334958 3556
rect 338666 3544 338672 3556
rect 338724 3544 338730 3596
rect 349246 3544 349252 3596
rect 349304 3584 349310 3596
rect 354030 3584 354036 3596
rect 349304 3556 354036 3584
rect 349304 3544 349310 3556
rect 354030 3544 354036 3556
rect 354088 3544 354094 3596
rect 373534 3544 373540 3596
rect 373592 3584 373598 3596
rect 379974 3584 379980 3596
rect 373592 3556 379980 3584
rect 373592 3544 373598 3556
rect 379974 3544 379980 3556
rect 380032 3544 380038 3596
rect 382366 3544 382372 3596
rect 382424 3584 382430 3596
rect 389450 3584 389456 3596
rect 382424 3556 389456 3584
rect 382424 3544 382430 3556
rect 389450 3544 389456 3556
rect 389508 3544 389514 3596
rect 390094 3544 390100 3596
rect 390152 3584 390158 3596
rect 397730 3584 397736 3596
rect 390152 3556 397736 3584
rect 390152 3544 390158 3556
rect 397730 3544 397736 3556
rect 397788 3544 397794 3596
rect 402238 3544 402244 3596
rect 402296 3584 402302 3596
rect 410794 3584 410800 3596
rect 402296 3556 410800 3584
rect 402296 3544 402302 3556
rect 410794 3544 410800 3556
rect 410852 3544 410858 3596
rect 412174 3544 412180 3596
rect 412232 3584 412238 3596
rect 421374 3584 421380 3596
rect 412232 3556 421380 3584
rect 412232 3544 412238 3556
rect 421374 3544 421380 3556
rect 421432 3544 421438 3596
rect 17034 3476 17040 3528
rect 17092 3516 17098 3528
rect 34606 3516 34612 3528
rect 17092 3488 34612 3516
rect 17092 3476 17098 3488
rect 34606 3476 34612 3488
rect 34664 3476 34670 3528
rect 45462 3476 45468 3528
rect 45520 3516 45526 3528
rect 61102 3516 61108 3528
rect 45520 3488 61108 3516
rect 45520 3476 45526 3488
rect 61102 3476 61108 3488
rect 61160 3476 61166 3528
rect 67910 3476 67916 3528
rect 67968 3516 67974 3528
rect 81710 3516 81716 3528
rect 67968 3488 81716 3516
rect 67968 3476 67974 3488
rect 81710 3476 81716 3488
rect 81768 3476 81774 3528
rect 86862 3476 86868 3528
rect 86920 3516 86926 3528
rect 99742 3516 99748 3528
rect 86920 3488 99748 3516
rect 86920 3476 86926 3488
rect 99742 3476 99748 3488
rect 99800 3476 99806 3528
rect 105722 3476 105728 3528
rect 105780 3516 105786 3528
rect 117406 3516 117412 3528
rect 105780 3488 117412 3516
rect 105780 3476 105786 3488
rect 117406 3476 117412 3488
rect 117464 3476 117470 3528
rect 129366 3476 129372 3528
rect 129424 3516 129430 3528
rect 139486 3516 139492 3528
rect 129424 3488 139492 3516
rect 129424 3476 129430 3488
rect 139486 3476 139492 3488
rect 139544 3476 139550 3528
rect 141234 3476 141240 3528
rect 141292 3516 141298 3528
rect 150526 3516 150532 3528
rect 141292 3488 150532 3516
rect 141292 3476 141298 3488
rect 150526 3476 150532 3488
rect 150584 3476 150590 3528
rect 153010 3476 153016 3528
rect 153068 3516 153074 3528
rect 161566 3516 161572 3528
rect 153068 3488 161572 3516
rect 153068 3476 153074 3488
rect 161566 3476 161572 3488
rect 161624 3476 161630 3528
rect 163682 3476 163688 3528
rect 163740 3516 163746 3528
rect 171502 3516 171508 3528
rect 163740 3488 171508 3516
rect 163740 3476 163746 3488
rect 171502 3476 171508 3488
rect 171560 3476 171566 3528
rect 187326 3476 187332 3528
rect 187384 3516 187390 3528
rect 193582 3516 193588 3528
rect 187384 3488 193588 3516
rect 187384 3476 187390 3488
rect 193582 3476 193588 3488
rect 193640 3476 193646 3528
rect 219250 3476 219256 3528
rect 219308 3516 219314 3528
rect 223390 3516 223396 3528
rect 219308 3488 223396 3516
rect 219308 3476 219314 3488
rect 223390 3476 223396 3488
rect 223448 3476 223454 3528
rect 372430 3476 372436 3528
rect 372488 3516 372494 3528
rect 378870 3516 378876 3528
rect 372488 3488 378876 3516
rect 372488 3476 372494 3488
rect 378870 3476 378876 3488
rect 378928 3476 378934 3528
rect 388990 3476 388996 3528
rect 389048 3516 389054 3528
rect 396534 3516 396540 3528
rect 389048 3488 396540 3516
rect 389048 3476 389054 3488
rect 396534 3476 396540 3488
rect 396592 3476 396598 3528
rect 404446 3476 404452 3528
rect 404504 3516 404510 3528
rect 413094 3516 413100 3528
rect 404504 3488 413100 3516
rect 404504 3476 404510 3488
rect 413094 3476 413100 3488
rect 413152 3476 413158 3528
rect 419902 3476 419908 3528
rect 419960 3516 419966 3528
rect 421852 3516 421880 3624
rect 429654 3612 429660 3624
rect 429712 3612 429718 3664
rect 443086 3612 443092 3664
rect 443144 3652 443150 3664
rect 454494 3652 454500 3664
rect 443144 3624 454500 3652
rect 443144 3612 443150 3624
rect 454494 3612 454500 3624
rect 454552 3612 454558 3664
rect 456334 3612 456340 3664
rect 456392 3652 456398 3664
rect 468294 3652 468300 3664
rect 456392 3624 468300 3652
rect 456392 3612 456398 3624
rect 468294 3612 468300 3624
rect 468352 3612 468358 3664
rect 468478 3612 468484 3664
rect 468536 3652 468542 3664
rect 481726 3652 481732 3664
rect 468536 3624 481732 3652
rect 468536 3612 468542 3624
rect 481726 3612 481732 3624
rect 481784 3612 481790 3664
rect 483934 3612 483940 3664
rect 483992 3652 483998 3664
rect 498194 3652 498200 3664
rect 483992 3624 498200 3652
rect 483992 3612 483998 3624
rect 498194 3612 498200 3624
rect 498252 3612 498258 3664
rect 499390 3612 499396 3664
rect 499448 3652 499454 3664
rect 514754 3652 514760 3664
rect 499448 3624 514760 3652
rect 499448 3612 499454 3624
rect 514754 3612 514760 3624
rect 514812 3612 514818 3664
rect 519262 3612 519268 3664
rect 519320 3652 519326 3664
rect 519320 3624 535776 3652
rect 519320 3612 519326 3624
rect 422110 3544 422116 3596
rect 422168 3584 422174 3596
rect 432046 3584 432052 3596
rect 422168 3556 432052 3584
rect 422168 3544 422174 3556
rect 432046 3544 432052 3556
rect 432104 3544 432110 3596
rect 433150 3544 433156 3596
rect 433208 3584 433214 3596
rect 443822 3584 443828 3596
rect 433208 3556 443828 3584
rect 433208 3544 433214 3556
rect 443822 3544 443828 3556
rect 443880 3544 443886 3596
rect 444190 3544 444196 3596
rect 444248 3584 444254 3596
rect 455690 3584 455696 3596
rect 444248 3556 455696 3584
rect 444248 3544 444254 3556
rect 455690 3544 455696 3556
rect 455748 3544 455754 3596
rect 465166 3584 465172 3596
rect 456996 3556 465172 3584
rect 422570 3516 422576 3528
rect 419960 3488 421880 3516
rect 422036 3488 422576 3516
rect 419960 3476 419966 3488
rect 4062 3408 4068 3460
rect 4120 3448 4126 3460
rect 22462 3448 22468 3460
rect 4120 3420 22468 3448
rect 4120 3408 4126 3420
rect 22462 3408 22468 3420
rect 22520 3408 22526 3460
rect 30098 3408 30104 3460
rect 30156 3448 30162 3460
rect 46750 3448 46756 3460
rect 30156 3420 46756 3448
rect 30156 3408 30162 3420
rect 46750 3408 46756 3420
rect 46808 3408 46814 3460
rect 48958 3408 48964 3460
rect 49016 3448 49022 3460
rect 64414 3448 64420 3460
rect 49016 3420 64420 3448
rect 49016 3408 49022 3420
rect 64414 3408 64420 3420
rect 64472 3408 64478 3460
rect 70302 3408 70308 3460
rect 70360 3448 70366 3460
rect 84286 3448 84292 3460
rect 70360 3420 84292 3448
rect 70360 3408 70366 3420
rect 84286 3408 84292 3420
rect 84344 3408 84350 3460
rect 87966 3408 87972 3460
rect 88024 3448 88030 3460
rect 100846 3448 100852 3460
rect 88024 3420 100852 3448
rect 88024 3408 88030 3420
rect 100846 3408 100852 3420
rect 100904 3408 100910 3460
rect 104526 3408 104532 3460
rect 104584 3448 104590 3460
rect 116302 3448 116308 3460
rect 104584 3420 116308 3448
rect 104584 3408 104590 3420
rect 116302 3408 116308 3420
rect 116360 3408 116366 3460
rect 121086 3408 121092 3460
rect 121144 3448 121150 3460
rect 131390 3448 131396 3460
rect 121144 3420 131396 3448
rect 121144 3408 121150 3420
rect 131390 3408 131396 3420
rect 131448 3408 131454 3460
rect 135254 3408 135260 3460
rect 135312 3448 135318 3460
rect 145006 3448 145012 3460
rect 135312 3420 145012 3448
rect 135312 3408 135318 3420
rect 145006 3408 145012 3420
rect 145064 3408 145070 3460
rect 147122 3408 147128 3460
rect 147180 3448 147186 3460
rect 156046 3448 156052 3460
rect 147180 3420 156052 3448
rect 147180 3408 147186 3420
rect 156046 3408 156052 3420
rect 156104 3408 156110 3460
rect 158898 3408 158904 3460
rect 158956 3448 158962 3460
rect 167086 3448 167092 3460
rect 158956 3420 167092 3448
rect 158956 3408 158962 3420
rect 167086 3408 167092 3420
rect 167144 3408 167150 3460
rect 170766 3408 170772 3460
rect 170824 3448 170830 3460
rect 178126 3448 178132 3460
rect 170824 3420 178132 3448
rect 170824 3408 170830 3420
rect 178126 3408 178132 3420
rect 178184 3408 178190 3460
rect 188522 3408 188528 3460
rect 188580 3448 188586 3460
rect 194686 3448 194692 3460
rect 188580 3420 194692 3448
rect 188580 3408 188586 3420
rect 194686 3408 194692 3420
rect 194744 3408 194750 3460
rect 199102 3408 199108 3460
rect 199160 3448 199166 3460
rect 204622 3448 204628 3460
rect 199160 3420 204628 3448
rect 199160 3408 199166 3420
rect 204622 3408 204628 3420
rect 204680 3408 204686 3460
rect 344830 3408 344836 3460
rect 344888 3448 344894 3460
rect 349246 3448 349252 3460
rect 344888 3420 349252 3448
rect 344888 3408 344894 3420
rect 349246 3408 349252 3420
rect 349304 3408 349310 3460
rect 352558 3408 352564 3460
rect 352616 3448 352622 3460
rect 357526 3448 357532 3460
rect 352616 3420 357532 3448
rect 352616 3408 352622 3420
rect 357526 3408 357532 3420
rect 357584 3408 357590 3460
rect 362494 3408 362500 3460
rect 362552 3448 362558 3460
rect 368198 3448 368204 3460
rect 362552 3420 368204 3448
rect 362552 3408 362558 3420
rect 368198 3408 368204 3420
rect 368256 3408 368262 3460
rect 383470 3408 383476 3460
rect 383528 3448 383534 3460
rect 390646 3448 390652 3460
rect 383528 3420 390652 3448
rect 383528 3408 383534 3420
rect 390646 3408 390652 3420
rect 390704 3408 390710 3460
rect 395614 3408 395620 3460
rect 395672 3448 395678 3460
rect 403618 3448 403624 3460
rect 395672 3420 403624 3448
rect 395672 3408 395678 3420
rect 403618 3408 403624 3420
rect 403676 3408 403682 3460
rect 406654 3408 406660 3460
rect 406712 3448 406718 3460
rect 415486 3448 415492 3460
rect 406712 3420 415492 3448
rect 406712 3408 406718 3420
rect 415486 3408 415492 3420
rect 415544 3408 415550 3460
rect 7650 3340 7656 3392
rect 7708 3380 7714 3392
rect 25774 3380 25780 3392
rect 7708 3352 25780 3380
rect 7708 3340 7714 3352
rect 25774 3340 25780 3352
rect 25832 3340 25838 3392
rect 33594 3340 33600 3392
rect 33652 3380 33658 3392
rect 50062 3380 50068 3392
rect 33652 3352 50068 3380
rect 33652 3340 33658 3352
rect 50062 3340 50068 3352
rect 50120 3340 50126 3392
rect 51350 3340 51356 3392
rect 51408 3380 51414 3392
rect 66622 3380 66628 3392
rect 51408 3352 66628 3380
rect 51408 3340 51414 3352
rect 66622 3340 66628 3352
rect 66680 3340 66686 3392
rect 76190 3340 76196 3392
rect 76248 3380 76254 3392
rect 89806 3380 89812 3392
rect 76248 3352 89812 3380
rect 76248 3340 76254 3352
rect 89806 3340 89812 3352
rect 89864 3340 89870 3392
rect 95142 3340 95148 3392
rect 95200 3380 95206 3392
rect 107470 3380 107476 3392
rect 95200 3352 107476 3380
rect 95200 3340 95206 3352
rect 107470 3340 107476 3352
rect 107528 3340 107534 3392
rect 118786 3340 118792 3392
rect 118844 3380 118850 3392
rect 129550 3380 129556 3392
rect 118844 3352 129556 3380
rect 118844 3340 118850 3352
rect 129550 3340 129556 3352
rect 129608 3340 129614 3392
rect 130562 3340 130568 3392
rect 130620 3380 130626 3392
rect 140590 3380 140596 3392
rect 130620 3352 140596 3380
rect 130620 3340 130626 3352
rect 140590 3340 140596 3352
rect 140648 3340 140654 3392
rect 392302 3340 392308 3392
rect 392360 3380 392366 3392
rect 400122 3380 400128 3392
rect 392360 3352 400128 3380
rect 392360 3340 392366 3352
rect 400122 3340 400128 3352
rect 400180 3340 400186 3392
rect 413278 3340 413284 3392
rect 413336 3380 413342 3392
rect 422036 3380 422064 3488
rect 422570 3476 422576 3488
rect 422628 3476 422634 3528
rect 428734 3476 428740 3528
rect 428792 3516 428798 3528
rect 439130 3516 439136 3528
rect 428792 3488 439136 3516
rect 428792 3476 428798 3488
rect 439130 3476 439136 3488
rect 439188 3476 439194 3528
rect 439774 3476 439780 3528
rect 439832 3516 439838 3528
rect 450906 3516 450912 3528
rect 439832 3488 450912 3516
rect 439832 3476 439838 3488
rect 450906 3476 450912 3488
rect 450964 3476 450970 3528
rect 453022 3476 453028 3528
rect 453080 3516 453086 3528
rect 456996 3516 457024 3556
rect 465166 3544 465172 3556
rect 465224 3544 465230 3596
rect 466270 3544 466276 3596
rect 466328 3584 466334 3596
rect 466328 3556 475240 3584
rect 466328 3544 466334 3556
rect 453080 3488 457024 3516
rect 453080 3476 453086 3488
rect 460750 3476 460756 3528
rect 460808 3516 460814 3528
rect 473446 3516 473452 3528
rect 460808 3488 473452 3516
rect 460808 3476 460814 3488
rect 473446 3476 473452 3488
rect 473504 3476 473510 3528
rect 428458 3448 428464 3460
rect 413336 3352 422064 3380
rect 422266 3420 428464 3448
rect 413336 3340 413342 3352
rect 2866 3272 2872 3324
rect 2924 3312 2930 3324
rect 21358 3312 21364 3324
rect 2924 3284 21364 3312
rect 2924 3272 2930 3284
rect 21358 3272 21364 3284
rect 21416 3272 21422 3324
rect 26510 3272 26516 3324
rect 26568 3312 26574 3324
rect 43438 3312 43444 3324
rect 26568 3284 43444 3312
rect 26568 3272 26574 3284
rect 43438 3272 43444 3284
rect 43496 3272 43502 3324
rect 53374 3312 53380 3324
rect 45526 3284 53380 3312
rect 12342 3204 12348 3256
rect 12400 3244 12406 3256
rect 30190 3244 30196 3256
rect 12400 3216 30196 3244
rect 12400 3204 12406 3216
rect 30190 3204 30196 3216
rect 30248 3204 30254 3256
rect 37182 3204 37188 3256
rect 37240 3244 37246 3256
rect 45526 3244 45554 3284
rect 53374 3272 53380 3284
rect 53432 3272 53438 3324
rect 54938 3272 54944 3324
rect 54996 3312 55002 3324
rect 69934 3312 69940 3324
rect 54996 3284 69940 3312
rect 54996 3272 55002 3284
rect 69934 3272 69940 3284
rect 69992 3272 69998 3324
rect 73798 3272 73804 3324
rect 73856 3312 73862 3324
rect 87598 3312 87604 3324
rect 73856 3284 87604 3312
rect 73856 3272 73862 3284
rect 87598 3272 87604 3284
rect 87656 3272 87662 3324
rect 109310 3272 109316 3324
rect 109368 3312 109374 3324
rect 120718 3312 120724 3324
rect 109368 3284 120724 3312
rect 109368 3272 109374 3284
rect 120718 3272 120724 3284
rect 120776 3272 120782 3324
rect 125870 3272 125876 3324
rect 125928 3312 125934 3324
rect 136174 3312 136180 3324
rect 125928 3284 136180 3312
rect 125928 3272 125934 3284
rect 136174 3272 136180 3284
rect 136232 3272 136238 3324
rect 365806 3272 365812 3324
rect 365864 3312 365870 3324
rect 371694 3312 371700 3324
rect 365864 3284 371700 3312
rect 365864 3272 365870 3284
rect 371694 3272 371700 3284
rect 371752 3272 371758 3324
rect 418798 3272 418804 3324
rect 418856 3312 418862 3324
rect 422266 3312 422294 3420
rect 428458 3408 428464 3420
rect 428516 3408 428522 3460
rect 429838 3408 429844 3460
rect 429896 3448 429902 3460
rect 440326 3448 440332 3460
rect 429896 3420 440332 3448
rect 429896 3408 429902 3420
rect 440326 3408 440332 3420
rect 440384 3408 440390 3460
rect 445294 3408 445300 3460
rect 445352 3448 445358 3460
rect 456886 3448 456892 3460
rect 445352 3420 456892 3448
rect 445352 3408 445358 3420
rect 456886 3408 456892 3420
rect 456944 3408 456950 3460
rect 459646 3408 459652 3460
rect 459704 3448 459710 3460
rect 472250 3448 472256 3460
rect 459704 3420 472256 3448
rect 459704 3408 459710 3420
rect 472250 3408 472256 3420
rect 472308 3408 472314 3460
rect 475212 3448 475240 3556
rect 479518 3544 479524 3596
rect 479576 3584 479582 3596
rect 493502 3584 493508 3596
rect 479576 3556 493508 3584
rect 479576 3544 479582 3556
rect 493502 3544 493508 3556
rect 493560 3544 493566 3596
rect 496078 3544 496084 3596
rect 496136 3584 496142 3596
rect 511258 3584 511264 3596
rect 496136 3556 511264 3584
rect 496136 3544 496142 3556
rect 511258 3544 511264 3556
rect 511316 3544 511322 3596
rect 512638 3544 512644 3596
rect 512696 3584 512702 3596
rect 529014 3584 529020 3596
rect 512696 3556 529020 3584
rect 512696 3544 512702 3556
rect 529014 3544 529020 3556
rect 529072 3544 529078 3596
rect 535748 3584 535776 3624
rect 535822 3612 535828 3664
rect 535880 3652 535886 3664
rect 553762 3652 553768 3664
rect 535880 3624 553768 3652
rect 535880 3612 535886 3624
rect 553762 3612 553768 3624
rect 553820 3612 553826 3664
rect 559006 3612 559012 3664
rect 559064 3652 559070 3664
rect 578602 3652 578608 3664
rect 559064 3624 578608 3652
rect 559064 3612 559070 3624
rect 578602 3612 578608 3624
rect 578660 3612 578666 3664
rect 536098 3584 536104 3596
rect 535748 3556 536104 3584
rect 536098 3544 536104 3556
rect 536156 3544 536162 3596
rect 543550 3544 543556 3596
rect 543608 3584 543614 3596
rect 562042 3584 562048 3596
rect 543608 3556 562048 3584
rect 543608 3544 543614 3556
rect 562042 3544 562048 3556
rect 562100 3544 562106 3596
rect 562318 3544 562324 3596
rect 562376 3584 562382 3596
rect 582190 3584 582196 3596
rect 562376 3556 582196 3584
rect 562376 3544 562382 3556
rect 582190 3544 582196 3556
rect 582248 3544 582254 3596
rect 475378 3476 475384 3528
rect 475436 3516 475442 3528
rect 480530 3516 480536 3528
rect 475436 3488 480536 3516
rect 475436 3476 475442 3488
rect 480530 3476 480536 3488
rect 480588 3476 480594 3528
rect 481634 3476 481640 3528
rect 481692 3516 481698 3528
rect 489914 3516 489920 3528
rect 481692 3488 489920 3516
rect 481692 3476 481698 3488
rect 489914 3476 489920 3488
rect 489972 3476 489978 3528
rect 490558 3476 490564 3528
rect 490616 3516 490622 3528
rect 505370 3516 505376 3528
rect 490616 3488 505376 3516
rect 490616 3476 490622 3488
rect 505370 3476 505376 3488
rect 505428 3476 505434 3528
rect 507118 3476 507124 3528
rect 507176 3516 507182 3528
rect 523034 3516 523040 3528
rect 507176 3488 523040 3516
rect 507176 3476 507182 3488
rect 523034 3476 523040 3488
rect 523092 3476 523098 3528
rect 523678 3476 523684 3528
rect 523736 3516 523742 3528
rect 526714 3516 526720 3528
rect 523736 3488 526720 3516
rect 523736 3476 523742 3488
rect 526714 3476 526720 3488
rect 526772 3476 526778 3528
rect 526990 3476 526996 3528
rect 527048 3516 527054 3528
rect 544378 3516 544384 3528
rect 527048 3488 544384 3516
rect 527048 3476 527054 3488
rect 544378 3476 544384 3488
rect 544436 3476 544442 3528
rect 544654 3476 544660 3528
rect 544712 3516 544718 3528
rect 563238 3516 563244 3528
rect 544712 3488 563244 3516
rect 544712 3476 544718 3488
rect 563238 3476 563244 3488
rect 563296 3476 563302 3528
rect 563422 3476 563428 3528
rect 563480 3516 563486 3528
rect 583386 3516 583392 3528
rect 563480 3488 583392 3516
rect 563480 3476 563486 3488
rect 583386 3476 583392 3488
rect 583444 3476 583450 3528
rect 479334 3448 479340 3460
rect 475212 3420 479340 3448
rect 479334 3408 479340 3420
rect 479392 3408 479398 3460
rect 486418 3448 486424 3460
rect 479444 3420 486424 3448
rect 438670 3340 438676 3392
rect 438728 3380 438734 3392
rect 449802 3380 449808 3392
rect 438728 3352 449808 3380
rect 438728 3340 438734 3352
rect 449802 3340 449808 3352
rect 449860 3340 449866 3392
rect 455230 3340 455236 3392
rect 455288 3380 455294 3392
rect 467466 3380 467472 3392
rect 455288 3352 467472 3380
rect 455288 3340 455294 3352
rect 467466 3340 467472 3352
rect 467524 3340 467530 3392
rect 469582 3340 469588 3392
rect 469640 3380 469646 3392
rect 469640 3352 470594 3380
rect 469640 3340 469646 3352
rect 418856 3284 422294 3312
rect 418856 3272 418862 3284
rect 447502 3272 447508 3324
rect 447560 3312 447566 3324
rect 459186 3312 459192 3324
rect 447560 3284 459192 3312
rect 447560 3272 447566 3284
rect 459186 3272 459192 3284
rect 459244 3272 459250 3324
rect 37240 3216 45554 3244
rect 37240 3204 37246 3216
rect 52546 3204 52552 3256
rect 52604 3244 52610 3256
rect 67726 3244 67732 3256
rect 52604 3216 67732 3244
rect 52604 3204 52610 3216
rect 67726 3204 67732 3216
rect 67784 3204 67790 3256
rect 72602 3204 72608 3256
rect 72660 3244 72666 3256
rect 86494 3244 86500 3256
rect 72660 3216 86500 3244
rect 72660 3204 72666 3216
rect 86494 3204 86500 3216
rect 86552 3204 86558 3256
rect 90358 3204 90364 3256
rect 90416 3244 90422 3256
rect 103054 3244 103060 3256
rect 90416 3216 103060 3244
rect 90416 3204 90422 3216
rect 103054 3204 103060 3216
rect 103112 3204 103118 3256
rect 106918 3204 106924 3256
rect 106976 3244 106982 3256
rect 118510 3244 118516 3256
rect 106976 3216 118516 3244
rect 106976 3204 106982 3216
rect 118510 3204 118516 3216
rect 118568 3204 118574 3256
rect 181438 3204 181444 3256
rect 181496 3244 181502 3256
rect 188062 3244 188068 3256
rect 181496 3216 188068 3244
rect 181496 3204 181502 3216
rect 188062 3204 188068 3216
rect 188120 3204 188126 3256
rect 201494 3204 201500 3256
rect 201552 3244 201558 3256
rect 206830 3244 206836 3256
rect 201552 3216 206836 3244
rect 201552 3204 201558 3216
rect 206830 3204 206836 3216
rect 206888 3204 206894 3256
rect 210970 3204 210976 3256
rect 211028 3244 211034 3256
rect 215662 3244 215668 3256
rect 211028 3216 215668 3244
rect 211028 3204 211034 3216
rect 215662 3204 215668 3216
rect 215720 3204 215726 3256
rect 331582 3204 331588 3256
rect 331640 3244 331646 3256
rect 335078 3244 335084 3256
rect 331640 3216 335084 3244
rect 331640 3204 331646 3216
rect 335078 3204 335084 3216
rect 335136 3204 335142 3256
rect 356974 3204 356980 3256
rect 357032 3244 357038 3256
rect 362310 3244 362316 3256
rect 357032 3216 362316 3244
rect 357032 3204 357038 3216
rect 362310 3204 362316 3216
rect 362368 3204 362374 3256
rect 440878 3204 440884 3256
rect 440936 3244 440942 3256
rect 452102 3244 452108 3256
rect 440936 3216 452108 3244
rect 440936 3204 440942 3216
rect 452102 3204 452108 3216
rect 452160 3204 452166 3256
rect 454126 3204 454132 3256
rect 454184 3244 454190 3256
rect 466270 3244 466276 3256
rect 454184 3216 466276 3244
rect 454184 3204 454190 3216
rect 466270 3204 466276 3216
rect 466328 3204 466334 3256
rect 24210 3136 24216 3188
rect 24268 3176 24274 3188
rect 41230 3176 41236 3188
rect 24268 3148 41236 3176
rect 24268 3136 24274 3148
rect 41230 3136 41236 3148
rect 41288 3136 41294 3188
rect 47854 3136 47860 3188
rect 47912 3176 47918 3188
rect 63310 3176 63316 3188
rect 47912 3148 63316 3176
rect 47912 3136 47918 3148
rect 63310 3136 63316 3148
rect 63368 3136 63374 3188
rect 65518 3136 65524 3188
rect 65576 3176 65582 3188
rect 79870 3176 79876 3188
rect 65576 3148 79876 3176
rect 65576 3136 65582 3148
rect 79870 3136 79876 3148
rect 79928 3136 79934 3188
rect 85666 3136 85672 3188
rect 85724 3176 85730 3188
rect 98270 3176 98276 3188
rect 85724 3148 98276 3176
rect 85724 3136 85730 3148
rect 98270 3136 98276 3148
rect 98328 3136 98334 3188
rect 182542 3136 182548 3188
rect 182600 3176 182606 3188
rect 189166 3176 189172 3188
rect 182600 3148 189172 3176
rect 182600 3136 182606 3148
rect 189166 3136 189172 3148
rect 189224 3136 189230 3188
rect 192018 3136 192024 3188
rect 192076 3176 192082 3188
rect 197998 3176 198004 3188
rect 192076 3148 198004 3176
rect 192076 3136 192082 3148
rect 197998 3136 198004 3148
rect 198056 3136 198062 3188
rect 203886 3136 203892 3188
rect 203944 3176 203950 3188
rect 209038 3176 209044 3188
rect 203944 3148 209044 3176
rect 203944 3136 203950 3148
rect 209038 3136 209044 3148
rect 209096 3136 209102 3188
rect 213362 3136 213368 3188
rect 213420 3176 213426 3188
rect 217870 3176 217876 3188
rect 213420 3148 217876 3176
rect 213420 3136 213426 3148
rect 217870 3136 217876 3148
rect 217928 3136 217934 3188
rect 223942 3136 223948 3188
rect 224000 3176 224006 3188
rect 227806 3176 227812 3188
rect 224000 3148 227812 3176
rect 224000 3136 224006 3148
rect 227806 3136 227812 3148
rect 227864 3136 227870 3188
rect 229830 3136 229836 3188
rect 229888 3176 229894 3188
rect 233326 3176 233332 3188
rect 229888 3148 233332 3176
rect 229888 3136 229894 3148
rect 233326 3136 233332 3148
rect 233384 3136 233390 3188
rect 246390 3136 246396 3188
rect 246448 3176 246454 3188
rect 248782 3176 248788 3188
rect 246448 3148 248788 3176
rect 246448 3136 246454 3148
rect 248782 3136 248788 3148
rect 248840 3136 248846 3188
rect 298462 3136 298468 3188
rect 298520 3176 298526 3188
rect 299658 3176 299664 3188
rect 298520 3148 299664 3176
rect 298520 3136 298526 3148
rect 299658 3136 299664 3148
rect 299716 3136 299722 3188
rect 322750 3136 322756 3188
rect 322808 3176 322814 3188
rect 325602 3176 325608 3188
rect 322808 3148 325608 3176
rect 322808 3136 322814 3148
rect 325602 3136 325608 3148
rect 325660 3136 325666 3188
rect 341518 3136 341524 3188
rect 341576 3176 341582 3188
rect 345750 3176 345756 3188
rect 341576 3148 345756 3176
rect 341576 3136 341582 3148
rect 345750 3136 345756 3148
rect 345808 3136 345814 3188
rect 348142 3136 348148 3188
rect 348200 3176 348206 3188
rect 352834 3176 352840 3188
rect 348200 3148 352840 3176
rect 348200 3136 348206 3148
rect 352834 3136 352840 3148
rect 352892 3136 352898 3188
rect 360286 3136 360292 3188
rect 360344 3176 360350 3188
rect 365806 3176 365812 3188
rect 360344 3148 365812 3176
rect 360344 3136 360350 3148
rect 365806 3136 365812 3148
rect 365864 3136 365870 3188
rect 370222 3136 370228 3188
rect 370280 3176 370286 3188
rect 376478 3176 376484 3188
rect 370280 3148 376484 3176
rect 370280 3136 370286 3148
rect 376478 3136 376484 3148
rect 376536 3136 376542 3188
rect 376846 3136 376852 3188
rect 376904 3176 376910 3188
rect 383562 3176 383568 3188
rect 376904 3148 383568 3176
rect 376904 3136 376910 3148
rect 383562 3136 383568 3148
rect 383620 3136 383626 3188
rect 384574 3136 384580 3188
rect 384632 3176 384638 3188
rect 391842 3176 391848 3188
rect 384632 3148 391848 3176
rect 384632 3136 384638 3148
rect 391842 3136 391848 3148
rect 391900 3136 391906 3188
rect 393406 3136 393412 3188
rect 393464 3176 393470 3188
rect 401318 3176 401324 3188
rect 393464 3148 401324 3176
rect 393464 3136 393470 3148
rect 401318 3136 401324 3148
rect 401376 3136 401382 3188
rect 449710 3136 449716 3188
rect 449768 3176 449774 3188
rect 461578 3176 461584 3188
rect 449768 3148 461584 3176
rect 449768 3136 449774 3148
rect 461578 3136 461584 3148
rect 461636 3136 461642 3188
rect 470566 3176 470594 3352
rect 472894 3272 472900 3324
rect 472952 3312 472958 3324
rect 479444 3312 479472 3420
rect 486418 3408 486424 3420
rect 486476 3408 486482 3460
rect 489454 3408 489460 3460
rect 489512 3448 489518 3460
rect 504174 3448 504180 3460
rect 489512 3420 504180 3448
rect 489512 3408 489518 3420
rect 504174 3408 504180 3420
rect 504232 3408 504238 3460
rect 506014 3408 506020 3460
rect 506072 3448 506078 3460
rect 521838 3448 521844 3460
rect 506072 3420 521844 3448
rect 506072 3408 506078 3420
rect 521838 3408 521844 3420
rect 521896 3408 521902 3460
rect 522574 3408 522580 3460
rect 522632 3448 522638 3460
rect 539594 3448 539600 3460
rect 522632 3420 539600 3448
rect 522632 3408 522638 3420
rect 539594 3408 539600 3420
rect 539652 3408 539658 3460
rect 542446 3408 542452 3460
rect 542504 3448 542510 3460
rect 560846 3448 560852 3460
rect 542504 3420 560852 3448
rect 542504 3408 542510 3420
rect 560846 3408 560852 3420
rect 560904 3408 560910 3460
rect 561214 3408 561220 3460
rect 561272 3448 561278 3460
rect 580994 3448 581000 3460
rect 561272 3420 581000 3448
rect 561272 3408 561278 3420
rect 580994 3408 581000 3420
rect 581052 3408 581058 3460
rect 482830 3380 482836 3392
rect 472952 3284 479472 3312
rect 479628 3352 482836 3380
rect 472952 3272 472958 3284
rect 479628 3176 479656 3352
rect 482830 3340 482836 3352
rect 482888 3340 482894 3392
rect 486142 3340 486148 3392
rect 486200 3380 486206 3392
rect 500586 3380 500592 3392
rect 486200 3352 500592 3380
rect 486200 3340 486206 3352
rect 500586 3340 500592 3352
rect 500644 3340 500650 3392
rect 500770 3340 500776 3392
rect 500828 3380 500834 3392
rect 515950 3380 515956 3392
rect 500828 3352 515956 3380
rect 500828 3340 500834 3352
rect 515950 3340 515956 3352
rect 516008 3340 516014 3392
rect 516042 3340 516048 3392
rect 516100 3380 516106 3392
rect 532510 3380 532516 3392
rect 516100 3352 532516 3380
rect 516100 3340 516106 3352
rect 532510 3340 532516 3352
rect 532568 3340 532574 3392
rect 532602 3340 532608 3392
rect 532660 3380 532666 3392
rect 550266 3380 550272 3392
rect 532660 3352 550272 3380
rect 532660 3340 532666 3352
rect 550266 3340 550272 3352
rect 550324 3340 550330 3392
rect 554590 3340 554596 3392
rect 554648 3380 554654 3392
rect 573910 3380 573916 3392
rect 554648 3352 573916 3380
rect 554648 3340 554654 3352
rect 573910 3340 573916 3352
rect 573968 3340 573974 3392
rect 484026 3312 484032 3324
rect 470566 3148 479656 3176
rect 480226 3284 484032 3312
rect 19426 3068 19432 3120
rect 19484 3108 19490 3120
rect 36814 3108 36820 3120
rect 19484 3080 36820 3108
rect 19484 3068 19490 3080
rect 36814 3068 36820 3080
rect 36872 3068 36878 3120
rect 44266 3068 44272 3120
rect 44324 3108 44330 3120
rect 59998 3108 60004 3120
rect 44324 3080 60004 3108
rect 44324 3068 44330 3080
rect 59998 3068 60004 3080
rect 60056 3068 60062 3120
rect 60826 3068 60832 3120
rect 60884 3108 60890 3120
rect 75454 3108 75460 3120
rect 60884 3080 75460 3108
rect 60884 3068 60890 3080
rect 75454 3068 75460 3080
rect 75512 3068 75518 3120
rect 102226 3068 102232 3120
rect 102284 3108 102290 3120
rect 114094 3108 114100 3120
rect 102284 3080 114100 3108
rect 102284 3068 102290 3080
rect 114094 3068 114100 3080
rect 114152 3068 114158 3120
rect 164878 3068 164884 3120
rect 164936 3108 164942 3120
rect 172606 3108 172612 3120
rect 164936 3080 172612 3108
rect 164936 3068 164942 3080
rect 172606 3068 172612 3080
rect 172664 3068 172670 3120
rect 184934 3068 184940 3120
rect 184992 3108 184998 3120
rect 191374 3108 191380 3120
rect 184992 3080 191380 3108
rect 184992 3068 184998 3080
rect 191374 3068 191380 3080
rect 191432 3068 191438 3120
rect 195606 3068 195612 3120
rect 195664 3108 195670 3120
rect 201310 3108 201316 3120
rect 195664 3080 201316 3108
rect 195664 3068 195670 3080
rect 201310 3068 201316 3080
rect 201368 3068 201374 3120
rect 205082 3068 205088 3120
rect 205140 3108 205146 3120
rect 210142 3108 210148 3120
rect 205140 3080 210148 3108
rect 205140 3068 205146 3080
rect 210142 3068 210148 3080
rect 210200 3068 210206 3120
rect 215662 3068 215668 3120
rect 215720 3108 215726 3120
rect 220078 3108 220084 3120
rect 215720 3080 220084 3108
rect 215720 3068 215726 3080
rect 220078 3068 220084 3080
rect 220136 3068 220142 3120
rect 221550 3068 221556 3120
rect 221608 3108 221614 3120
rect 225598 3108 225604 3120
rect 221608 3080 225604 3108
rect 221608 3068 221614 3080
rect 225598 3068 225604 3080
rect 225656 3068 225662 3120
rect 226334 3068 226340 3120
rect 226392 3108 226398 3120
rect 230014 3108 230020 3120
rect 226392 3080 230020 3108
rect 226392 3068 226398 3080
rect 230014 3068 230020 3080
rect 230072 3068 230078 3120
rect 231026 3068 231032 3120
rect 231084 3108 231090 3120
rect 234430 3108 234436 3120
rect 231084 3080 234436 3108
rect 231084 3068 231090 3080
rect 234430 3068 234436 3080
rect 234488 3068 234494 3120
rect 234614 3068 234620 3120
rect 234672 3108 234678 3120
rect 237742 3108 237748 3120
rect 234672 3080 237748 3108
rect 234672 3068 234678 3080
rect 237742 3068 237748 3080
rect 237800 3068 237806 3120
rect 238110 3068 238116 3120
rect 238168 3108 238174 3120
rect 241054 3108 241060 3120
rect 238168 3080 241060 3108
rect 238168 3068 238174 3080
rect 241054 3068 241060 3080
rect 241112 3068 241118 3120
rect 241698 3068 241704 3120
rect 241756 3108 241762 3120
rect 244366 3108 244372 3120
rect 241756 3080 244372 3108
rect 241756 3068 241762 3080
rect 244366 3068 244372 3080
rect 244424 3068 244430 3120
rect 247586 3068 247592 3120
rect 247644 3108 247650 3120
rect 249886 3108 249892 3120
rect 247644 3080 249892 3108
rect 247644 3068 247650 3080
rect 249886 3068 249892 3080
rect 249944 3068 249950 3120
rect 249978 3068 249984 3120
rect 250036 3108 250042 3120
rect 252094 3108 252100 3120
rect 250036 3080 252100 3108
rect 250036 3068 250042 3080
rect 252094 3068 252100 3080
rect 252152 3068 252158 3120
rect 252370 3068 252376 3120
rect 252428 3108 252434 3120
rect 254302 3108 254308 3120
rect 252428 3080 254308 3108
rect 252428 3068 252434 3080
rect 254302 3068 254308 3080
rect 254360 3068 254366 3120
rect 254670 3068 254676 3120
rect 254728 3108 254734 3120
rect 256510 3108 256516 3120
rect 254728 3080 256516 3108
rect 254728 3068 254734 3080
rect 256510 3068 256516 3080
rect 256568 3068 256574 3120
rect 257062 3068 257068 3120
rect 257120 3108 257126 3120
rect 258718 3108 258724 3120
rect 257120 3080 258724 3108
rect 257120 3068 257126 3080
rect 258718 3068 258724 3080
rect 258776 3068 258782 3120
rect 259454 3068 259460 3120
rect 259512 3108 259518 3120
rect 260926 3108 260932 3120
rect 259512 3080 260932 3108
rect 259512 3068 259518 3080
rect 260926 3068 260932 3080
rect 260984 3068 260990 3120
rect 261754 3068 261760 3120
rect 261812 3108 261818 3120
rect 263134 3108 263140 3120
rect 261812 3080 263140 3108
rect 261812 3068 261818 3080
rect 263134 3068 263140 3080
rect 263192 3068 263198 3120
rect 264146 3068 264152 3120
rect 264204 3108 264210 3120
rect 265342 3108 265348 3120
rect 264204 3080 265348 3108
rect 264204 3068 264210 3080
rect 265342 3068 265348 3080
rect 265400 3068 265406 3120
rect 271230 3068 271236 3120
rect 271288 3108 271294 3120
rect 271966 3108 271972 3120
rect 271288 3080 271972 3108
rect 271288 3068 271294 3080
rect 271966 3068 271972 3080
rect 272024 3068 272030 3120
rect 300670 3068 300676 3120
rect 300728 3108 300734 3120
rect 301958 3108 301964 3120
rect 300728 3080 301964 3108
rect 300728 3068 300734 3080
rect 301958 3068 301964 3080
rect 302016 3068 302022 3120
rect 302878 3068 302884 3120
rect 302936 3108 302942 3120
rect 304350 3108 304356 3120
rect 302936 3080 304356 3108
rect 302936 3068 302942 3080
rect 304350 3068 304356 3080
rect 304408 3068 304414 3120
rect 305086 3068 305092 3120
rect 305144 3108 305150 3120
rect 306742 3108 306748 3120
rect 305144 3080 306748 3108
rect 305144 3068 305150 3080
rect 306742 3068 306748 3080
rect 306800 3068 306806 3120
rect 307294 3068 307300 3120
rect 307352 3108 307358 3120
rect 309042 3108 309048 3120
rect 307352 3080 309048 3108
rect 307352 3068 307358 3080
rect 309042 3068 309048 3080
rect 309100 3068 309106 3120
rect 311710 3068 311716 3120
rect 311768 3108 311774 3120
rect 313826 3108 313832 3120
rect 311768 3080 313832 3108
rect 311768 3068 311774 3080
rect 313826 3068 313832 3080
rect 313884 3068 313890 3120
rect 315022 3068 315028 3120
rect 315080 3108 315086 3120
rect 317322 3108 317328 3120
rect 315080 3080 317328 3108
rect 315080 3068 315086 3080
rect 317322 3068 317328 3080
rect 317380 3068 317386 3120
rect 319438 3068 319444 3120
rect 319496 3108 319502 3120
rect 322106 3108 322112 3120
rect 319496 3080 322112 3108
rect 319496 3068 319502 3080
rect 322106 3068 322112 3080
rect 322164 3068 322170 3120
rect 324958 3068 324964 3120
rect 325016 3108 325022 3120
rect 327994 3108 328000 3120
rect 325016 3080 328000 3108
rect 325016 3068 325022 3080
rect 327994 3068 328000 3080
rect 328052 3068 328058 3120
rect 328270 3068 328276 3120
rect 328328 3108 328334 3120
rect 331582 3108 331588 3120
rect 328328 3080 331588 3108
rect 328328 3068 328334 3080
rect 331582 3068 331588 3080
rect 331640 3068 331646 3120
rect 332686 3068 332692 3120
rect 332744 3108 332750 3120
rect 336274 3108 336280 3120
rect 332744 3080 336280 3108
rect 332744 3068 332750 3080
rect 336274 3068 336280 3080
rect 336332 3068 336338 3120
rect 337102 3068 337108 3120
rect 337160 3108 337166 3120
rect 340966 3108 340972 3120
rect 337160 3080 340972 3108
rect 337160 3068 337166 3080
rect 340966 3068 340972 3080
rect 341024 3068 341030 3120
rect 345934 3068 345940 3120
rect 345992 3108 345998 3120
rect 350442 3108 350448 3120
rect 345992 3080 350448 3108
rect 345992 3068 345998 3080
rect 350442 3068 350448 3080
rect 350500 3068 350506 3120
rect 359182 3068 359188 3120
rect 359240 3108 359246 3120
rect 364610 3108 364616 3120
rect 359240 3080 364616 3108
rect 359240 3068 359246 3080
rect 364610 3068 364616 3080
rect 364668 3068 364674 3120
rect 369118 3068 369124 3120
rect 369176 3108 369182 3120
rect 375282 3108 375288 3120
rect 369176 3080 375288 3108
rect 369176 3068 369182 3080
rect 375282 3068 375288 3080
rect 375340 3068 375346 3120
rect 379054 3068 379060 3120
rect 379112 3108 379118 3120
rect 385954 3108 385960 3120
rect 379112 3080 385960 3108
rect 379112 3068 379118 3080
rect 385954 3068 385960 3080
rect 386012 3068 386018 3120
rect 386782 3068 386788 3120
rect 386840 3108 386846 3120
rect 394234 3108 394240 3120
rect 386840 3080 394240 3108
rect 386840 3068 386846 3080
rect 394234 3068 394240 3080
rect 394292 3068 394298 3120
rect 403342 3068 403348 3120
rect 403400 3108 403406 3120
rect 411898 3108 411904 3120
rect 403400 3080 411904 3108
rect 403400 3068 403406 3080
rect 411898 3068 411904 3080
rect 411956 3068 411962 3120
rect 470686 3068 470692 3120
rect 470744 3108 470750 3120
rect 480226 3108 480254 3284
rect 484026 3272 484032 3284
rect 484084 3272 484090 3324
rect 487246 3272 487252 3324
rect 487304 3312 487310 3324
rect 501782 3312 501788 3324
rect 487304 3284 501788 3312
rect 487304 3272 487310 3284
rect 501782 3272 501788 3284
rect 501840 3272 501846 3324
rect 501874 3272 501880 3324
rect 501932 3312 501938 3324
rect 517146 3312 517152 3324
rect 501932 3284 517152 3312
rect 501932 3272 501938 3284
rect 517146 3272 517152 3284
rect 517204 3272 517210 3324
rect 524782 3272 524788 3324
rect 524840 3312 524846 3324
rect 524840 3284 526668 3312
rect 524840 3272 524846 3284
rect 492766 3204 492772 3256
rect 492824 3244 492830 3256
rect 507670 3244 507676 3256
rect 492824 3216 507676 3244
rect 492824 3204 492830 3216
rect 507670 3204 507676 3216
rect 507728 3204 507734 3256
rect 509326 3204 509332 3256
rect 509384 3244 509390 3256
rect 525426 3244 525432 3256
rect 509384 3216 525432 3244
rect 509384 3204 509390 3216
rect 525426 3204 525432 3216
rect 525484 3204 525490 3256
rect 526640 3244 526668 3284
rect 526714 3272 526720 3324
rect 526772 3312 526778 3324
rect 540790 3312 540796 3324
rect 526772 3284 540796 3312
rect 526772 3272 526778 3284
rect 540790 3272 540796 3284
rect 540848 3272 540854 3324
rect 558546 3312 558552 3324
rect 544028 3284 558552 3312
rect 541986 3244 541992 3256
rect 526640 3216 541992 3244
rect 541986 3204 541992 3216
rect 542044 3204 542050 3256
rect 485038 3136 485044 3188
rect 485096 3176 485102 3188
rect 499390 3176 499396 3188
rect 485096 3148 499396 3176
rect 485096 3136 485102 3148
rect 499390 3136 499396 3148
rect 499448 3136 499454 3188
rect 517054 3136 517060 3188
rect 517112 3176 517118 3188
rect 533706 3176 533712 3188
rect 517112 3148 533712 3176
rect 517112 3136 517118 3148
rect 533706 3136 533712 3148
rect 533764 3136 533770 3188
rect 540238 3136 540244 3188
rect 540296 3176 540302 3188
rect 544028 3176 544056 3284
rect 558546 3272 558552 3284
rect 558604 3272 558610 3324
rect 546862 3204 546868 3256
rect 546920 3244 546926 3256
rect 565630 3244 565636 3256
rect 546920 3216 565636 3244
rect 546920 3204 546926 3216
rect 565630 3204 565636 3216
rect 565688 3204 565694 3256
rect 559742 3176 559748 3188
rect 540296 3148 544056 3176
rect 552676 3148 559748 3176
rect 540296 3136 540302 3148
rect 470744 3080 480254 3108
rect 470744 3068 470750 3080
rect 480622 3068 480628 3120
rect 480680 3108 480686 3120
rect 494698 3108 494704 3120
rect 480680 3080 494704 3108
rect 480680 3068 480686 3080
rect 494698 3068 494704 3080
rect 494756 3068 494762 3120
rect 503806 3068 503812 3120
rect 503864 3108 503870 3120
rect 519538 3108 519544 3120
rect 503864 3080 519544 3108
rect 503864 3068 503870 3080
rect 519538 3068 519544 3080
rect 519596 3068 519602 3120
rect 531406 3068 531412 3120
rect 531464 3108 531470 3120
rect 549070 3108 549076 3120
rect 531464 3080 549076 3108
rect 531464 3068 531470 3080
rect 549070 3068 549076 3080
rect 549128 3068 549134 3120
rect 18230 3000 18236 3052
rect 18288 3040 18294 3052
rect 35710 3040 35716 3052
rect 18288 3012 35716 3040
rect 18288 3000 18294 3012
rect 35710 3000 35716 3012
rect 35768 3000 35774 3052
rect 69106 3000 69112 3052
rect 69164 3040 69170 3052
rect 83182 3040 83188 3052
rect 69164 3012 83188 3040
rect 69164 3000 69170 3012
rect 83182 3000 83188 3012
rect 83240 3000 83246 3052
rect 142430 3000 142436 3052
rect 142488 3040 142494 3052
rect 151630 3040 151636 3052
rect 142488 3012 151636 3040
rect 142488 3000 142494 3012
rect 151630 3000 151636 3012
rect 151688 3000 151694 3052
rect 151814 3000 151820 3052
rect 151872 3040 151878 3052
rect 160462 3040 160468 3052
rect 151872 3012 160468 3040
rect 151872 3000 151878 3012
rect 160462 3000 160468 3012
rect 160520 3000 160526 3052
rect 166074 3000 166080 3052
rect 166132 3040 166138 3052
rect 173710 3040 173716 3052
rect 166132 3012 173716 3040
rect 166132 3000 166138 3012
rect 173710 3000 173716 3012
rect 173768 3000 173774 3052
rect 186130 3000 186136 3052
rect 186188 3040 186194 3052
rect 192478 3040 192484 3052
rect 186188 3012 192484 3040
rect 186188 3000 186194 3012
rect 192478 3000 192484 3012
rect 192536 3000 192542 3052
rect 196802 3000 196808 3052
rect 196860 3040 196866 3052
rect 202414 3040 202420 3052
rect 196860 3012 202420 3040
rect 196860 3000 196866 3012
rect 202414 3000 202420 3012
rect 202472 3000 202478 3052
rect 207382 3000 207388 3052
rect 207440 3040 207446 3052
rect 212350 3040 212356 3052
rect 207440 3012 212356 3040
rect 207440 3000 207446 3012
rect 212350 3000 212356 3012
rect 212408 3000 212414 3052
rect 216858 3000 216864 3052
rect 216916 3040 216922 3052
rect 221182 3040 221188 3052
rect 216916 3012 221188 3040
rect 216916 3000 216922 3012
rect 221182 3000 221188 3012
rect 221240 3000 221246 3052
rect 222746 3000 222752 3052
rect 222804 3040 222810 3052
rect 226702 3040 226708 3052
rect 222804 3012 226708 3040
rect 222804 3000 222810 3012
rect 226702 3000 226708 3012
rect 226760 3000 226766 3052
rect 227530 3000 227536 3052
rect 227588 3040 227594 3052
rect 231118 3040 231124 3052
rect 227588 3012 231124 3040
rect 227588 3000 227594 3012
rect 231118 3000 231124 3012
rect 231176 3000 231182 3052
rect 233418 3000 233424 3052
rect 233476 3040 233482 3052
rect 236638 3040 236644 3052
rect 233476 3012 236644 3040
rect 233476 3000 233482 3012
rect 236638 3000 236644 3012
rect 236696 3000 236702 3052
rect 237006 3000 237012 3052
rect 237064 3040 237070 3052
rect 239950 3040 239956 3052
rect 237064 3012 239956 3040
rect 237064 3000 237070 3012
rect 239950 3000 239956 3012
rect 240008 3000 240014 3052
rect 240502 3000 240508 3052
rect 240560 3040 240566 3052
rect 243262 3040 243268 3052
rect 240560 3012 243268 3040
rect 240560 3000 240566 3012
rect 243262 3000 243268 3012
rect 243320 3000 243326 3052
rect 244090 3000 244096 3052
rect 244148 3040 244154 3052
rect 246574 3040 246580 3052
rect 244148 3012 246580 3040
rect 244148 3000 244154 3012
rect 246574 3000 246580 3012
rect 246632 3000 246638 3052
rect 248782 3000 248788 3052
rect 248840 3040 248846 3052
rect 250990 3040 250996 3052
rect 248840 3012 250996 3040
rect 248840 3000 248846 3012
rect 250990 3000 250996 3012
rect 251048 3000 251054 3052
rect 251174 3000 251180 3052
rect 251232 3040 251238 3052
rect 253198 3040 253204 3052
rect 251232 3012 253204 3040
rect 251232 3000 251238 3012
rect 253198 3000 253204 3012
rect 253256 3000 253262 3052
rect 253474 3000 253480 3052
rect 253532 3040 253538 3052
rect 255406 3040 255412 3052
rect 253532 3012 255412 3040
rect 253532 3000 253538 3012
rect 255406 3000 255412 3012
rect 255464 3000 255470 3052
rect 255866 3000 255872 3052
rect 255924 3040 255930 3052
rect 257614 3040 257620 3052
rect 255924 3012 257620 3040
rect 255924 3000 255930 3012
rect 257614 3000 257620 3012
rect 257672 3000 257678 3052
rect 258258 3000 258264 3052
rect 258316 3040 258322 3052
rect 259822 3040 259828 3052
rect 258316 3012 259828 3040
rect 258316 3000 258322 3012
rect 259822 3000 259828 3012
rect 259880 3000 259886 3052
rect 260650 3000 260656 3052
rect 260708 3040 260714 3052
rect 262030 3040 262036 3052
rect 260708 3012 262036 3040
rect 260708 3000 260714 3012
rect 262030 3000 262036 3012
rect 262088 3000 262094 3052
rect 262950 3000 262956 3052
rect 263008 3040 263014 3052
rect 264238 3040 264244 3052
rect 263008 3012 264244 3040
rect 263008 3000 263014 3012
rect 264238 3000 264244 3012
rect 264296 3000 264302 3052
rect 267734 3000 267740 3052
rect 267792 3040 267798 3052
rect 268654 3040 268660 3052
rect 267792 3012 268660 3040
rect 267792 3000 267798 3012
rect 268654 3000 268660 3012
rect 268712 3000 268718 3052
rect 291838 3000 291844 3052
rect 291896 3040 291902 3052
rect 292574 3040 292580 3052
rect 291896 3012 292580 3040
rect 291896 3000 291902 3012
rect 292574 3000 292580 3012
rect 292632 3000 292638 3052
rect 294046 3000 294052 3052
rect 294104 3040 294110 3052
rect 294874 3040 294880 3052
rect 294104 3012 294880 3040
rect 294104 3000 294110 3012
rect 294874 3000 294880 3012
rect 294932 3000 294938 3052
rect 295150 3000 295156 3052
rect 295208 3040 295214 3052
rect 296070 3040 296076 3052
rect 295208 3012 296076 3040
rect 295208 3000 295214 3012
rect 296070 3000 296076 3012
rect 296128 3000 296134 3052
rect 296254 3000 296260 3052
rect 296312 3040 296318 3052
rect 297266 3040 297272 3052
rect 296312 3012 297272 3040
rect 296312 3000 296318 3012
rect 297266 3000 297272 3012
rect 297324 3000 297330 3052
rect 297358 3000 297364 3052
rect 297416 3040 297422 3052
rect 298462 3040 298468 3052
rect 297416 3012 298468 3040
rect 297416 3000 297422 3012
rect 298462 3000 298468 3012
rect 298520 3000 298526 3052
rect 299566 3000 299572 3052
rect 299624 3040 299630 3052
rect 300762 3040 300768 3052
rect 299624 3012 300768 3040
rect 299624 3000 299630 3012
rect 300762 3000 300768 3012
rect 300820 3000 300826 3052
rect 301774 3000 301780 3052
rect 301832 3040 301838 3052
rect 303154 3040 303160 3052
rect 301832 3012 303160 3040
rect 301832 3000 301838 3012
rect 303154 3000 303160 3012
rect 303212 3000 303218 3052
rect 303982 3000 303988 3052
rect 304040 3040 304046 3052
rect 305546 3040 305552 3052
rect 304040 3012 305552 3040
rect 304040 3000 304046 3012
rect 305546 3000 305552 3012
rect 305604 3000 305610 3052
rect 306190 3000 306196 3052
rect 306248 3040 306254 3052
rect 307938 3040 307944 3052
rect 306248 3012 307944 3040
rect 306248 3000 306254 3012
rect 307938 3000 307944 3012
rect 307996 3000 308002 3052
rect 308398 3000 308404 3052
rect 308456 3040 308462 3052
rect 310238 3040 310244 3052
rect 308456 3012 310244 3040
rect 308456 3000 308462 3012
rect 310238 3000 310244 3012
rect 310296 3000 310302 3052
rect 310606 3000 310612 3052
rect 310664 3040 310670 3052
rect 312630 3040 312636 3052
rect 310664 3012 312636 3040
rect 310664 3000 310670 3012
rect 312630 3000 312636 3012
rect 312688 3000 312694 3052
rect 313918 3000 313924 3052
rect 313976 3040 313982 3052
rect 316218 3040 316224 3052
rect 313976 3012 316224 3040
rect 313976 3000 313982 3012
rect 316218 3000 316224 3012
rect 316276 3000 316282 3052
rect 317230 3000 317236 3052
rect 317288 3040 317294 3052
rect 319714 3040 319720 3052
rect 317288 3012 319720 3040
rect 317288 3000 317294 3012
rect 319714 3000 319720 3012
rect 319772 3000 319778 3052
rect 320542 3000 320548 3052
rect 320600 3040 320606 3052
rect 323302 3040 323308 3052
rect 320600 3012 323308 3040
rect 320600 3000 320606 3012
rect 323302 3000 323308 3012
rect 323360 3000 323366 3052
rect 326062 3000 326068 3052
rect 326120 3040 326126 3052
rect 329190 3040 329196 3052
rect 326120 3012 329196 3040
rect 326120 3000 326126 3012
rect 329190 3000 329196 3012
rect 329248 3000 329254 3052
rect 330478 3000 330484 3052
rect 330536 3040 330542 3052
rect 333882 3040 333888 3052
rect 330536 3012 333888 3040
rect 330536 3000 330542 3012
rect 333882 3000 333888 3012
rect 333940 3000 333946 3052
rect 335998 3000 336004 3052
rect 336056 3040 336062 3052
rect 339862 3040 339868 3052
rect 336056 3012 339868 3040
rect 336056 3000 336062 3012
rect 339862 3000 339868 3012
rect 339920 3000 339926 3052
rect 340414 3000 340420 3052
rect 340472 3040 340478 3052
rect 344554 3040 344560 3052
rect 340472 3012 344560 3040
rect 340472 3000 340478 3012
rect 344554 3000 344560 3012
rect 344612 3000 344618 3052
rect 347038 3000 347044 3052
rect 347096 3040 347102 3052
rect 351638 3040 351644 3052
rect 347096 3012 351644 3040
rect 347096 3000 347102 3012
rect 351638 3000 351644 3012
rect 351696 3000 351702 3052
rect 354766 3000 354772 3052
rect 354824 3040 354830 3052
rect 359918 3040 359924 3052
rect 354824 3012 359924 3040
rect 354824 3000 354830 3012
rect 359918 3000 359924 3012
rect 359976 3000 359982 3052
rect 364702 3000 364708 3052
rect 364760 3040 364766 3052
rect 370590 3040 370596 3052
rect 364760 3012 370596 3040
rect 364760 3000 364766 3012
rect 370590 3000 370596 3012
rect 370648 3000 370654 3052
rect 374638 3000 374644 3052
rect 374696 3040 374702 3052
rect 381170 3040 381176 3052
rect 374696 3012 381176 3040
rect 374696 3000 374702 3012
rect 381170 3000 381176 3012
rect 381228 3000 381234 3052
rect 387886 3000 387892 3052
rect 387944 3040 387950 3052
rect 395338 3040 395344 3052
rect 387944 3012 395344 3040
rect 387944 3000 387950 3012
rect 395338 3000 395344 3012
rect 395396 3000 395402 3052
rect 396718 3000 396724 3052
rect 396776 3040 396782 3052
rect 404814 3040 404820 3052
rect 396776 3012 404820 3040
rect 396776 3000 396782 3012
rect 404814 3000 404820 3012
rect 404872 3000 404878 3052
rect 508222 3000 508228 3052
rect 508280 3040 508286 3052
rect 524230 3040 524236 3052
rect 508280 3012 524236 3040
rect 508280 3000 508286 3012
rect 524230 3000 524236 3012
rect 524288 3000 524294 3052
rect 541342 3000 541348 3052
rect 541400 3040 541406 3052
rect 552676 3040 552704 3148
rect 559742 3136 559748 3148
rect 559800 3136 559806 3188
rect 566826 3108 566832 3120
rect 541400 3012 552704 3040
rect 557506 3080 566832 3108
rect 541400 3000 541406 3012
rect 25314 2932 25320 2984
rect 25372 2972 25378 2984
rect 42334 2972 42340 2984
rect 25372 2944 42340 2972
rect 25372 2932 25378 2944
rect 42334 2932 42340 2944
rect 42392 2932 42398 2984
rect 59630 2932 59636 2984
rect 59688 2972 59694 2984
rect 74350 2972 74356 2984
rect 59688 2944 74356 2972
rect 59688 2932 59694 2944
rect 74350 2932 74356 2944
rect 74408 2932 74414 2984
rect 162486 2932 162492 2984
rect 162544 2972 162550 2984
rect 170398 2972 170404 2984
rect 162544 2944 170404 2972
rect 162544 2932 162550 2944
rect 170398 2932 170404 2944
rect 170456 2932 170462 2984
rect 171962 2932 171968 2984
rect 172020 2972 172026 2984
rect 179230 2972 179236 2984
rect 172020 2944 179236 2972
rect 172020 2932 172026 2944
rect 179230 2932 179236 2944
rect 179288 2932 179294 2984
rect 183738 2932 183744 2984
rect 183796 2972 183802 2984
rect 190270 2972 190276 2984
rect 183796 2944 190276 2972
rect 183796 2932 183802 2944
rect 190270 2932 190276 2944
rect 190328 2932 190334 2984
rect 194410 2932 194416 2984
rect 194468 2972 194474 2984
rect 200206 2972 200212 2984
rect 194468 2944 200212 2972
rect 194468 2932 194474 2944
rect 200206 2932 200212 2944
rect 200264 2932 200270 2984
rect 200298 2932 200304 2984
rect 200356 2972 200362 2984
rect 205726 2972 205732 2984
rect 200356 2944 205732 2972
rect 200356 2932 200362 2944
rect 205726 2932 205732 2944
rect 205784 2932 205790 2984
rect 206186 2932 206192 2984
rect 206244 2972 206250 2984
rect 211246 2972 211252 2984
rect 206244 2944 211252 2972
rect 206244 2932 206250 2944
rect 211246 2932 211252 2944
rect 211304 2932 211310 2984
rect 214466 2932 214472 2984
rect 214524 2972 214530 2984
rect 218974 2972 218980 2984
rect 214524 2944 218980 2972
rect 214524 2932 214530 2944
rect 218974 2932 218980 2944
rect 219032 2932 219038 2984
rect 220446 2932 220452 2984
rect 220504 2972 220510 2984
rect 224494 2972 224500 2984
rect 220504 2944 224500 2972
rect 220504 2932 220510 2944
rect 224494 2932 224500 2944
rect 224552 2932 224558 2984
rect 225138 2932 225144 2984
rect 225196 2972 225202 2984
rect 228910 2972 228916 2984
rect 225196 2944 228916 2972
rect 225196 2932 225202 2944
rect 228910 2932 228916 2944
rect 228968 2932 228974 2984
rect 232222 2932 232228 2984
rect 232280 2972 232286 2984
rect 235534 2972 235540 2984
rect 232280 2944 235540 2972
rect 232280 2932 232286 2944
rect 235534 2932 235540 2944
rect 235592 2932 235598 2984
rect 239306 2932 239312 2984
rect 239364 2972 239370 2984
rect 242158 2972 242164 2984
rect 239364 2944 242164 2972
rect 239364 2932 239370 2944
rect 242158 2932 242164 2944
rect 242216 2932 242222 2984
rect 245194 2932 245200 2984
rect 245252 2972 245258 2984
rect 247678 2972 247684 2984
rect 245252 2944 247684 2972
rect 245252 2932 245258 2944
rect 247678 2932 247684 2944
rect 247736 2932 247742 2984
rect 316126 2932 316132 2984
rect 316184 2972 316190 2984
rect 318518 2972 318524 2984
rect 316184 2944 318524 2972
rect 316184 2932 316190 2944
rect 318518 2932 318524 2944
rect 318576 2932 318582 2984
rect 323854 2932 323860 2984
rect 323912 2972 323918 2984
rect 326798 2972 326804 2984
rect 323912 2944 326804 2972
rect 323912 2932 323918 2944
rect 326798 2932 326804 2944
rect 326856 2932 326862 2984
rect 327166 2932 327172 2984
rect 327224 2972 327230 2984
rect 330386 2972 330392 2984
rect 327224 2944 330392 2972
rect 327224 2932 327230 2944
rect 330386 2932 330392 2944
rect 330444 2932 330450 2984
rect 333790 2932 333796 2984
rect 333848 2972 333854 2984
rect 337470 2972 337476 2984
rect 333848 2944 337476 2972
rect 333848 2932 333854 2944
rect 337470 2932 337476 2944
rect 337528 2932 337534 2984
rect 338206 2932 338212 2984
rect 338264 2972 338270 2984
rect 342162 2972 342168 2984
rect 338264 2944 342168 2972
rect 338264 2932 338270 2944
rect 342162 2932 342168 2944
rect 342220 2932 342226 2984
rect 342622 2932 342628 2984
rect 342680 2972 342686 2984
rect 346946 2972 346952 2984
rect 342680 2944 346952 2972
rect 342680 2932 342686 2944
rect 346946 2932 346952 2944
rect 347004 2932 347010 2984
rect 351454 2932 351460 2984
rect 351512 2972 351518 2984
rect 356330 2972 356336 2984
rect 351512 2944 356336 2972
rect 351512 2932 351518 2944
rect 356330 2932 356336 2944
rect 356388 2932 356394 2984
rect 361390 2932 361396 2984
rect 361448 2972 361454 2984
rect 367002 2972 367008 2984
rect 361448 2944 367008 2972
rect 361448 2932 361454 2944
rect 367002 2932 367008 2944
rect 367060 2932 367066 2984
rect 368014 2932 368020 2984
rect 368072 2972 368078 2984
rect 374086 2972 374092 2984
rect 368072 2944 374092 2972
rect 368072 2932 368078 2944
rect 374086 2932 374092 2944
rect 374144 2932 374150 2984
rect 377950 2932 377956 2984
rect 378008 2972 378014 2984
rect 384758 2972 384764 2984
rect 378008 2944 384764 2972
rect 378008 2932 378014 2944
rect 384758 2932 384764 2944
rect 384816 2932 384822 2984
rect 385678 2932 385684 2984
rect 385736 2972 385742 2984
rect 393038 2972 393044 2984
rect 385736 2944 393044 2972
rect 385736 2932 385742 2944
rect 393038 2932 393044 2944
rect 393096 2932 393102 2984
rect 394510 2932 394516 2984
rect 394568 2972 394574 2984
rect 402514 2972 402520 2984
rect 394568 2944 402520 2972
rect 394568 2932 394574 2944
rect 402514 2932 402520 2944
rect 402572 2932 402578 2984
rect 547966 2932 547972 2984
rect 548024 2972 548030 2984
rect 557506 2972 557534 3080
rect 566826 3068 566832 3080
rect 566884 3068 566890 3120
rect 548024 2944 557534 2972
rect 548024 2932 548030 2944
rect 27706 2864 27712 2916
rect 27764 2904 27770 2916
rect 44542 2904 44548 2916
rect 27764 2876 44548 2904
rect 27764 2864 27770 2876
rect 44542 2864 44548 2876
rect 44600 2864 44606 2916
rect 155402 2864 155408 2916
rect 155460 2904 155466 2916
rect 163774 2904 163780 2916
rect 155460 2876 163780 2904
rect 155460 2864 155466 2876
rect 163774 2864 163780 2876
rect 163832 2864 163838 2916
rect 173158 2864 173164 2916
rect 173216 2904 173222 2916
rect 180334 2904 180340 2916
rect 173216 2876 180340 2904
rect 173216 2864 173222 2876
rect 180334 2864 180340 2876
rect 180392 2864 180398 2916
rect 190822 2864 190828 2916
rect 190880 2904 190886 2916
rect 196894 2904 196900 2916
rect 190880 2876 196900 2904
rect 190880 2864 190886 2876
rect 196894 2864 196900 2876
rect 196952 2864 196958 2916
rect 202690 2864 202696 2916
rect 202748 2904 202754 2916
rect 207934 2904 207940 2916
rect 202748 2876 207940 2904
rect 202748 2864 202754 2876
rect 207934 2864 207940 2876
rect 207992 2864 207998 2916
rect 212166 2864 212172 2916
rect 212224 2904 212230 2916
rect 216766 2904 216772 2916
rect 212224 2876 216772 2904
rect 212224 2864 212230 2876
rect 216766 2864 216772 2876
rect 216824 2864 216830 2916
rect 235810 2864 235816 2916
rect 235868 2904 235874 2916
rect 238846 2904 238852 2916
rect 235868 2876 238852 2904
rect 235868 2864 235874 2876
rect 238846 2864 238852 2876
rect 238904 2864 238910 2916
rect 242894 2864 242900 2916
rect 242952 2904 242958 2916
rect 245470 2904 245476 2916
rect 242952 2876 245476 2904
rect 242952 2864 242958 2876
rect 245470 2864 245476 2876
rect 245528 2864 245534 2916
rect 265342 2864 265348 2916
rect 265400 2904 265406 2916
rect 266446 2904 266452 2916
rect 265400 2876 266452 2904
rect 265400 2864 265406 2876
rect 266446 2864 266452 2876
rect 266504 2864 266510 2916
rect 268838 2864 268844 2916
rect 268896 2904 268902 2916
rect 269758 2904 269764 2916
rect 268896 2876 269764 2904
rect 268896 2864 268902 2876
rect 269758 2864 269764 2876
rect 269816 2864 269822 2916
rect 329374 2864 329380 2916
rect 329432 2904 329438 2916
rect 332686 2904 332692 2916
rect 329432 2876 332692 2904
rect 329432 2864 329438 2876
rect 332686 2864 332692 2876
rect 332744 2864 332750 2916
rect 339310 2864 339316 2916
rect 339368 2904 339374 2916
rect 343358 2904 343364 2916
rect 339368 2876 343364 2904
rect 339368 2864 339374 2876
rect 343358 2864 343364 2876
rect 343416 2864 343422 2916
rect 350350 2864 350356 2916
rect 350408 2904 350414 2916
rect 355226 2904 355232 2916
rect 350408 2876 355232 2904
rect 350408 2864 350414 2876
rect 355226 2864 355232 2876
rect 355284 2864 355290 2916
rect 355870 2864 355876 2916
rect 355928 2904 355934 2916
rect 361114 2904 361120 2916
rect 355928 2876 361120 2904
rect 355928 2864 355934 2876
rect 361114 2864 361120 2876
rect 361172 2864 361178 2916
rect 375742 2864 375748 2916
rect 375800 2904 375806 2916
rect 382366 2904 382372 2916
rect 375800 2876 382372 2904
rect 375800 2864 375806 2876
rect 382366 2864 382372 2876
rect 382424 2864 382430 2916
rect 35986 2796 35992 2848
rect 36044 2836 36050 2848
rect 52270 2836 52276 2848
rect 36044 2808 52276 2836
rect 36044 2796 36050 2808
rect 52270 2796 52276 2808
rect 52328 2796 52334 2848
rect 209774 2796 209780 2848
rect 209832 2836 209838 2848
rect 214558 2836 214564 2848
rect 209832 2808 214564 2836
rect 209832 2796 209838 2808
rect 214558 2796 214564 2808
rect 214616 2796 214622 2848
rect 309502 2796 309508 2848
rect 309560 2836 309566 2848
rect 311434 2836 311440 2848
rect 309560 2808 311440 2836
rect 309560 2796 309566 2808
rect 311434 2796 311440 2808
rect 311492 2796 311498 2848
rect 312814 2796 312820 2848
rect 312872 2836 312878 2848
rect 315022 2836 315028 2848
rect 312872 2808 315028 2836
rect 312872 2796 312878 2808
rect 315022 2796 315028 2808
rect 315080 2796 315086 2848
rect 318334 2796 318340 2848
rect 318392 2836 318398 2848
rect 320910 2836 320916 2848
rect 318392 2808 320916 2836
rect 318392 2796 318398 2808
rect 320910 2796 320916 2808
rect 320968 2796 320974 2848
rect 321646 2796 321652 2848
rect 321704 2836 321710 2848
rect 324406 2836 324412 2848
rect 321704 2808 324412 2836
rect 321704 2796 321710 2808
rect 324406 2796 324412 2808
rect 324464 2796 324470 2848
rect 358078 2796 358084 2848
rect 358136 2836 358142 2848
rect 363506 2836 363512 2848
rect 358136 2808 363512 2836
rect 358136 2796 358142 2808
rect 363506 2796 363512 2808
rect 363564 2796 363570 2848
rect 366910 2796 366916 2848
rect 366968 2836 366974 2848
rect 372890 2836 372896 2848
rect 366968 2808 372896 2836
rect 366968 2796 366974 2808
rect 372890 2796 372896 2808
rect 372948 2796 372954 2848
rect 474734 2796 474740 2848
rect 474792 2836 474798 2848
rect 475746 2836 475752 2848
rect 474792 2808 475752 2836
rect 474792 2796 474798 2808
rect 475746 2796 475752 2808
rect 475804 2796 475810 2848
rect 525794 2796 525800 2848
rect 525852 2836 525858 2848
rect 526622 2836 526628 2848
rect 525852 2808 526628 2836
rect 525852 2796 525858 2808
rect 526622 2796 526628 2808
rect 526680 2796 526686 2848
<< via1 >>
rect 201500 702992 201552 703044
rect 202788 702992 202840 703044
rect 105452 700884 105504 700936
rect 109040 700884 109092 700936
rect 89168 700680 89220 700732
rect 93032 700680 93084 700732
rect 56784 700476 56836 700528
rect 61384 700476 61436 700528
rect 40500 700340 40552 700392
rect 44180 700340 44232 700392
rect 8116 700272 8168 700324
rect 13912 700272 13964 700324
rect 24308 699660 24360 699712
rect 28264 699660 28316 699712
rect 72976 699660 73028 699712
rect 76104 699660 76156 699712
rect 137836 699660 137888 699712
rect 140780 699660 140832 699712
rect 298744 699660 298796 699712
rect 300124 699660 300176 699712
rect 314660 699660 314712 699712
rect 316316 699660 316368 699712
rect 330392 699660 330444 699712
rect 332508 699660 332560 699712
rect 346400 699660 346452 699712
rect 348792 699660 348844 699712
rect 362040 699660 362092 699712
rect 364984 699660 365036 699712
rect 378140 699660 378192 699712
rect 381176 699660 381228 699712
rect 393688 699660 393740 699712
rect 397460 699660 397512 699712
rect 409880 699660 409932 699712
rect 413652 699660 413704 699712
rect 425336 699660 425388 699712
rect 429844 699660 429896 699712
rect 441620 699660 441672 699712
rect 446128 699660 446180 699712
rect 574100 699660 574152 699712
rect 575848 699660 575900 699712
rect 28264 695444 28316 695496
rect 30196 695444 30248 695496
rect 76104 695444 76156 695496
rect 77668 695444 77720 695496
rect 153200 695444 153252 695496
rect 156788 695444 156840 695496
rect 186504 695444 186556 695496
rect 188436 695444 188488 695496
rect 201500 695444 201552 695496
rect 204260 695444 204312 695496
rect 520740 695444 520792 695496
rect 527180 695444 527232 695496
rect 473268 695376 473320 695428
rect 477500 695376 477552 695428
rect 568212 695240 568264 695292
rect 574100 695240 574152 695292
rect 489092 694764 489144 694816
rect 494060 694764 494112 694816
rect 536564 694764 536616 694816
rect 542360 694764 542412 694816
rect 44180 694152 44232 694204
rect 46020 694152 46072 694204
rect 121644 694152 121696 694204
rect 125140 694152 125192 694204
rect 169760 694152 169812 694204
rect 172612 694152 172664 694204
rect 218060 694152 218112 694204
rect 220084 694152 220136 694204
rect 457444 694152 457496 694204
rect 462320 694152 462372 694204
rect 504916 694152 504968 694204
rect 510620 694152 510672 694204
rect 552388 694152 552440 694204
rect 558920 694152 558972 694204
rect 578332 672936 578384 672988
rect 580264 672936 580316 672988
rect 578516 659404 578568 659456
rect 580264 659404 580316 659456
rect 578332 646960 578384 647012
rect 580264 646960 580316 647012
rect 578332 620916 578384 620968
rect 580264 620916 580316 620968
rect 578240 510620 578292 510672
rect 580540 510620 580592 510672
rect 578240 470976 578292 471028
rect 579804 470976 579856 471028
rect 578240 404336 578292 404388
rect 580356 404336 580408 404388
rect 578332 362720 578384 362772
rect 580908 362720 580960 362772
rect 578516 219716 578568 219768
rect 580908 219716 580960 219768
rect 578332 181296 578384 181348
rect 580540 181296 580592 181348
rect 578792 142536 578844 142588
rect 580724 142536 580776 142588
rect 578332 116696 578384 116748
rect 580264 116696 580316 116748
rect 578240 60664 578292 60716
rect 580816 60664 580868 60716
rect 578240 20612 578292 20664
rect 580632 20612 580684 20664
rect 1676 4088 1728 4140
rect 20260 4088 20312 4140
rect 21824 4088 21876 4140
rect 39028 4088 39080 4140
rect 43076 4088 43128 4140
rect 58900 4088 58952 4140
rect 66720 4088 66772 4140
rect 80980 4088 81032 4140
rect 83280 4088 83332 4140
rect 96436 4088 96488 4140
rect 97448 4088 97500 4140
rect 109684 4088 109736 4140
rect 112812 4088 112864 4140
rect 124036 4088 124088 4140
rect 124680 4088 124732 4140
rect 135076 4088 135128 4140
rect 136456 4088 136508 4140
rect 146116 4088 146168 4140
rect 157800 4088 157852 4140
rect 165988 4088 166040 4140
rect 174268 4088 174320 4140
rect 181444 4088 181496 4140
rect 415492 4088 415544 4140
rect 424968 4088 425020 4140
rect 430948 4088 431000 4140
rect 441528 4088 441580 4140
rect 464068 4088 464120 4140
rect 476948 4088 477000 4140
rect 477316 4088 477368 4140
rect 491116 4088 491168 4140
rect 493876 4088 493928 4140
rect 508872 4088 508924 4140
rect 510436 4088 510488 4140
rect 525800 4088 525852 4140
rect 525892 4088 525944 4140
rect 543188 4088 543240 4140
rect 549076 4088 549128 4140
rect 568028 4088 568080 4140
rect 15936 4020 15988 4072
rect 33508 4020 33560 4072
rect 40684 4020 40736 4072
rect 56692 4020 56744 4072
rect 62028 4020 62080 4072
rect 76564 4020 76616 4072
rect 77392 4020 77444 4072
rect 90916 4020 90968 4072
rect 93952 4020 94004 4072
rect 106372 4020 106424 4072
rect 119896 4020 119948 4072
rect 130660 4020 130712 4072
rect 132960 4020 133012 4072
rect 142804 4020 142856 4072
rect 143540 4020 143592 4072
rect 152740 4020 152792 4072
rect 154212 4020 154264 4072
rect 162676 4020 162728 4072
rect 168380 4020 168432 4072
rect 175924 4020 175976 4072
rect 176660 4020 176712 4072
rect 183652 4020 183704 4072
rect 400036 4020 400088 4072
rect 408408 4020 408460 4072
rect 421012 4020 421064 4072
rect 430856 4020 430908 4072
rect 432052 4020 432104 4072
rect 442632 4020 442684 4072
rect 448612 4020 448664 4072
rect 460388 4020 460440 4072
rect 465172 4020 465224 4072
rect 6460 3952 6512 4004
rect 24676 3952 24728 4004
rect 39580 3952 39632 4004
rect 55588 3952 55640 4004
rect 58440 3952 58492 4004
rect 73252 3952 73304 4004
rect 84476 3952 84528 4004
rect 97540 3952 97592 4004
rect 101036 3952 101088 4004
rect 112996 3952 113048 4004
rect 115296 3952 115348 4004
rect 126244 3952 126296 4004
rect 126980 3952 127032 4004
rect 137284 3952 137336 4004
rect 150624 3952 150676 4004
rect 159364 3952 159416 4004
rect 180248 3952 180300 4004
rect 186964 3952 187016 4004
rect 189724 3952 189776 4004
rect 195796 3952 195848 4004
rect 407764 3952 407816 4004
rect 13544 3884 13596 3936
rect 31300 3884 31352 3936
rect 38384 3884 38436 3936
rect 54484 3884 54536 3936
rect 57244 3884 57296 3936
rect 72148 3884 72200 3936
rect 78588 3884 78640 3936
rect 92020 3884 92072 3936
rect 92756 3884 92808 3936
rect 105268 3884 105320 3936
rect 108120 3884 108172 3936
rect 119620 3884 119672 3936
rect 122288 3884 122340 3936
rect 132868 3884 132920 3936
rect 134156 3884 134208 3936
rect 143908 3884 143960 3936
rect 149520 3884 149572 3936
rect 158260 3884 158312 3936
rect 160100 3884 160152 3936
rect 168196 3884 168248 3936
rect 179052 3884 179104 3936
rect 185860 3884 185912 3936
rect 401140 3884 401192 3936
rect 8760 3816 8812 3868
rect 26884 3816 26936 3868
rect 32496 3816 32548 3868
rect 48964 3816 49016 3868
rect 53748 3816 53800 3868
rect 68836 3816 68888 3868
rect 71504 3816 71556 3868
rect 85396 3816 85448 3868
rect 89168 3816 89220 3868
rect 101956 3816 102008 3868
rect 103336 3816 103388 3868
rect 115204 3816 115256 3868
rect 116400 3816 116452 3868
rect 127348 3816 127400 3868
rect 137652 3816 137704 3868
rect 147220 3816 147272 3868
rect 148324 3816 148376 3868
rect 157156 3816 157208 3868
rect 161296 3816 161348 3868
rect 169300 3816 169352 3868
rect 353668 3816 353720 3868
rect 358728 3816 358780 3868
rect 371332 3816 371384 3868
rect 377680 3816 377732 3868
rect 397828 3816 397880 3868
rect 406016 3816 406068 3868
rect 408868 3884 408920 3936
rect 416596 3952 416648 4004
rect 426164 3952 426216 4004
rect 426532 3952 426584 4004
rect 436744 3952 436796 4004
rect 437572 3952 437624 4004
rect 448520 3952 448572 4004
rect 461860 3952 461912 4004
rect 474556 3952 474608 4004
rect 476212 4020 476264 4072
rect 481640 4020 481692 4072
rect 481732 4020 481784 4072
rect 495900 4020 495952 4072
rect 498292 4020 498344 4072
rect 513564 4020 513616 4072
rect 520372 4020 520424 4072
rect 536840 4020 536892 4072
rect 536932 4020 536984 4072
rect 554964 4020 555016 4072
rect 556804 4020 556856 4072
rect 576308 4020 576360 4072
rect 478144 3952 478196 4004
rect 478420 3952 478472 4004
rect 492312 3952 492364 4004
rect 497188 3952 497240 4004
rect 512460 3952 512512 4004
rect 513748 3952 513800 4004
rect 530124 3952 530176 4004
rect 530308 3952 530360 4004
rect 547880 3952 547932 4004
rect 550180 3952 550232 4004
rect 569132 3952 569184 4004
rect 409604 3816 409656 3868
rect 409972 3816 410024 3868
rect 416688 3884 416740 3936
rect 417700 3884 417752 3936
rect 427268 3884 427320 3936
rect 427636 3884 427688 3936
rect 437940 3884 437992 3936
rect 441988 3884 442040 3936
rect 453304 3884 453356 3936
rect 457444 3884 457496 3936
rect 469864 3884 469916 3936
rect 471796 3884 471848 3936
rect 485228 3884 485280 3936
rect 488356 3884 488408 3936
rect 572 3748 624 3800
rect 19156 3748 19208 3800
rect 23020 3748 23072 3800
rect 40132 3748 40184 3800
rect 41880 3748 41932 3800
rect 57796 3748 57848 3800
rect 63224 3748 63276 3800
rect 77668 3748 77720 3800
rect 79692 3748 79744 3800
rect 93124 3748 93176 3800
rect 96252 3748 96304 3800
rect 108580 3748 108632 3800
rect 110512 3748 110564 3800
rect 121828 3748 121880 3800
rect 123484 3748 123536 3800
rect 133972 3748 134024 3800
rect 140044 3748 140096 3800
rect 149428 3748 149480 3800
rect 167184 3748 167236 3800
rect 174820 3748 174872 3800
rect 175464 3748 175516 3800
rect 182548 3748 182600 3800
rect 197912 3748 197964 3800
rect 203524 3748 203576 3800
rect 208584 3748 208636 3800
rect 213460 3748 213512 3800
rect 218060 3748 218112 3800
rect 222292 3748 222344 3800
rect 381268 3748 381320 3800
rect 388260 3748 388312 3800
rect 398932 3748 398984 3800
rect 407212 3748 407264 3800
rect 411076 3748 411128 3800
rect 417884 3816 417936 3868
rect 424324 3816 424376 3868
rect 434444 3816 434496 3868
rect 434536 3816 434588 3868
rect 445024 3816 445076 3868
rect 446404 3816 446456 3868
rect 458088 3816 458140 3868
rect 458548 3816 458600 3868
rect 471060 3816 471112 3868
rect 474004 3816 474056 3868
rect 487620 3816 487672 3868
rect 9956 3680 10008 3732
rect 27988 3680 28040 3732
rect 31300 3680 31352 3732
rect 47860 3680 47912 3732
rect 50160 3680 50212 3732
rect 65524 3680 65576 3732
rect 75000 3680 75052 3732
rect 88708 3680 88760 3732
rect 91560 3680 91612 3732
rect 104164 3680 104216 3732
rect 117596 3680 117648 3732
rect 128452 3680 128504 3732
rect 138848 3680 138900 3732
rect 147956 3680 148008 3732
rect 177856 3680 177908 3732
rect 184756 3680 184808 3732
rect 228732 3680 228784 3732
rect 232228 3680 232280 3732
rect 418988 3748 419040 3800
rect 423220 3748 423272 3800
rect 433248 3748 433300 3800
rect 435364 3748 435416 3800
rect 446220 3748 446272 3800
rect 451924 3748 451976 3800
rect 463976 3748 464028 3800
rect 467380 3748 467432 3800
rect 475384 3748 475436 3800
rect 482836 3748 482888 3800
rect 497096 3816 497148 3868
rect 502708 3884 502760 3936
rect 517980 3884 518032 3936
rect 518164 3884 518216 3936
rect 534540 3884 534592 3936
rect 534724 3884 534776 3936
rect 552664 3884 552716 3936
rect 553492 3884 553544 3936
rect 572720 3884 572772 3936
rect 502984 3816 503036 3868
rect 491668 3748 491720 3800
rect 506480 3816 506532 3868
rect 514852 3816 514904 3868
rect 531320 3816 531372 3868
rect 533620 3816 533672 3868
rect 551100 3816 551152 3868
rect 551284 3816 551336 3868
rect 570328 3816 570380 3868
rect 504916 3748 504968 3800
rect 520740 3748 520792 3800
rect 529204 3748 529256 3800
rect 546684 3748 546736 3800
rect 557908 3748 557960 3800
rect 577412 3748 577464 3800
rect 420184 3680 420236 3732
rect 14740 3612 14792 3664
rect 32404 3612 32456 3664
rect 34796 3612 34848 3664
rect 51172 3612 51224 3664
rect 56048 3612 56100 3664
rect 71044 3612 71096 3664
rect 82084 3612 82136 3664
rect 95332 3612 95384 3664
rect 99840 3612 99892 3664
rect 111892 3612 111944 3664
rect 114008 3612 114060 3664
rect 125140 3612 125192 3664
rect 131764 3612 131816 3664
rect 141700 3612 141752 3664
rect 144736 3612 144788 3664
rect 153844 3612 153896 3664
rect 343732 3612 343784 3664
rect 348056 3612 348108 3664
rect 363604 3612 363656 3664
rect 369400 3612 369452 3664
rect 380164 3612 380216 3664
rect 387156 3612 387208 3664
rect 391204 3612 391256 3664
rect 398932 3612 398984 3664
rect 405556 3612 405608 3664
rect 414296 3612 414348 3664
rect 414388 3612 414440 3664
rect 423772 3680 423824 3732
rect 425428 3680 425480 3732
rect 435548 3680 435600 3732
rect 436468 3680 436520 3732
rect 447416 3680 447468 3732
rect 450820 3680 450872 3732
rect 462780 3680 462832 3732
rect 462964 3680 463016 3732
rect 474740 3680 474792 3732
rect 475476 3680 475528 3732
rect 488816 3680 488868 3732
rect 494980 3680 495032 3732
rect 510068 3680 510120 3732
rect 511540 3680 511592 3732
rect 527824 3680 527876 3732
rect 528100 3680 528152 3732
rect 545488 3680 545540 3732
rect 545764 3680 545816 3732
rect 564440 3680 564492 3732
rect 11152 3544 11204 3596
rect 29092 3544 29144 3596
rect 46664 3544 46716 3596
rect 62212 3544 62264 3596
rect 64328 3544 64380 3596
rect 78772 3544 78824 3596
rect 80888 3544 80940 3596
rect 94228 3544 94280 3596
rect 98644 3544 98696 3596
rect 110788 3544 110840 3596
rect 111616 3544 111668 3596
rect 122932 3544 122984 3596
rect 128176 3544 128228 3596
rect 138388 3544 138440 3596
rect 145932 3544 145984 3596
rect 154948 3544 155000 3596
rect 156604 3544 156656 3596
rect 164884 3544 164936 3596
rect 169576 3544 169628 3596
rect 177028 3544 177080 3596
rect 193220 3544 193272 3596
rect 199108 3544 199160 3596
rect 334900 3544 334952 3596
rect 338672 3544 338724 3596
rect 349252 3544 349304 3596
rect 354036 3544 354088 3596
rect 373540 3544 373592 3596
rect 379980 3544 380032 3596
rect 382372 3544 382424 3596
rect 389456 3544 389508 3596
rect 390100 3544 390152 3596
rect 397736 3544 397788 3596
rect 402244 3544 402296 3596
rect 410800 3544 410852 3596
rect 412180 3544 412232 3596
rect 421380 3544 421432 3596
rect 17040 3476 17092 3528
rect 34612 3476 34664 3528
rect 45468 3476 45520 3528
rect 61108 3476 61160 3528
rect 67916 3476 67968 3528
rect 81716 3476 81768 3528
rect 86868 3476 86920 3528
rect 99748 3476 99800 3528
rect 105728 3476 105780 3528
rect 117412 3476 117464 3528
rect 129372 3476 129424 3528
rect 139492 3476 139544 3528
rect 141240 3476 141292 3528
rect 150532 3476 150584 3528
rect 153016 3476 153068 3528
rect 161572 3476 161624 3528
rect 163688 3476 163740 3528
rect 171508 3476 171560 3528
rect 187332 3476 187384 3528
rect 193588 3476 193640 3528
rect 219256 3476 219308 3528
rect 223396 3476 223448 3528
rect 372436 3476 372488 3528
rect 378876 3476 378928 3528
rect 388996 3476 389048 3528
rect 396540 3476 396592 3528
rect 404452 3476 404504 3528
rect 413100 3476 413152 3528
rect 419908 3476 419960 3528
rect 429660 3612 429712 3664
rect 443092 3612 443144 3664
rect 454500 3612 454552 3664
rect 456340 3612 456392 3664
rect 468300 3612 468352 3664
rect 468484 3612 468536 3664
rect 481732 3612 481784 3664
rect 483940 3612 483992 3664
rect 498200 3612 498252 3664
rect 499396 3612 499448 3664
rect 514760 3612 514812 3664
rect 519268 3612 519320 3664
rect 422116 3544 422168 3596
rect 432052 3544 432104 3596
rect 433156 3544 433208 3596
rect 443828 3544 443880 3596
rect 444196 3544 444248 3596
rect 455696 3544 455748 3596
rect 4068 3408 4120 3460
rect 22468 3408 22520 3460
rect 30104 3408 30156 3460
rect 46756 3408 46808 3460
rect 48964 3408 49016 3460
rect 64420 3408 64472 3460
rect 70308 3408 70360 3460
rect 84292 3408 84344 3460
rect 87972 3408 88024 3460
rect 100852 3408 100904 3460
rect 104532 3408 104584 3460
rect 116308 3408 116360 3460
rect 121092 3408 121144 3460
rect 131396 3408 131448 3460
rect 135260 3408 135312 3460
rect 145012 3408 145064 3460
rect 147128 3408 147180 3460
rect 156052 3408 156104 3460
rect 158904 3408 158956 3460
rect 167092 3408 167144 3460
rect 170772 3408 170824 3460
rect 178132 3408 178184 3460
rect 188528 3408 188580 3460
rect 194692 3408 194744 3460
rect 199108 3408 199160 3460
rect 204628 3408 204680 3460
rect 344836 3408 344888 3460
rect 349252 3408 349304 3460
rect 352564 3408 352616 3460
rect 357532 3408 357584 3460
rect 362500 3408 362552 3460
rect 368204 3408 368256 3460
rect 383476 3408 383528 3460
rect 390652 3408 390704 3460
rect 395620 3408 395672 3460
rect 403624 3408 403676 3460
rect 406660 3408 406712 3460
rect 415492 3408 415544 3460
rect 7656 3340 7708 3392
rect 25780 3340 25832 3392
rect 33600 3340 33652 3392
rect 50068 3340 50120 3392
rect 51356 3340 51408 3392
rect 66628 3340 66680 3392
rect 76196 3340 76248 3392
rect 89812 3340 89864 3392
rect 95148 3340 95200 3392
rect 107476 3340 107528 3392
rect 118792 3340 118844 3392
rect 129556 3340 129608 3392
rect 130568 3340 130620 3392
rect 140596 3340 140648 3392
rect 392308 3340 392360 3392
rect 400128 3340 400180 3392
rect 413284 3340 413336 3392
rect 422576 3476 422628 3528
rect 428740 3476 428792 3528
rect 439136 3476 439188 3528
rect 439780 3476 439832 3528
rect 450912 3476 450964 3528
rect 453028 3476 453080 3528
rect 465172 3544 465224 3596
rect 466276 3544 466328 3596
rect 460756 3476 460808 3528
rect 473452 3476 473504 3528
rect 2872 3272 2924 3324
rect 21364 3272 21416 3324
rect 26516 3272 26568 3324
rect 43444 3272 43496 3324
rect 12348 3204 12400 3256
rect 30196 3204 30248 3256
rect 37188 3204 37240 3256
rect 53380 3272 53432 3324
rect 54944 3272 54996 3324
rect 69940 3272 69992 3324
rect 73804 3272 73856 3324
rect 87604 3272 87656 3324
rect 109316 3272 109368 3324
rect 120724 3272 120776 3324
rect 125876 3272 125928 3324
rect 136180 3272 136232 3324
rect 365812 3272 365864 3324
rect 371700 3272 371752 3324
rect 418804 3272 418856 3324
rect 428464 3408 428516 3460
rect 429844 3408 429896 3460
rect 440332 3408 440384 3460
rect 445300 3408 445352 3460
rect 456892 3408 456944 3460
rect 459652 3408 459704 3460
rect 472256 3408 472308 3460
rect 479524 3544 479576 3596
rect 493508 3544 493560 3596
rect 496084 3544 496136 3596
rect 511264 3544 511316 3596
rect 512644 3544 512696 3596
rect 529020 3544 529072 3596
rect 535828 3612 535880 3664
rect 553768 3612 553820 3664
rect 559012 3612 559064 3664
rect 578608 3612 578660 3664
rect 536104 3544 536156 3596
rect 543556 3544 543608 3596
rect 562048 3544 562100 3596
rect 562324 3544 562376 3596
rect 582196 3544 582248 3596
rect 475384 3476 475436 3528
rect 480536 3476 480588 3528
rect 481640 3476 481692 3528
rect 489920 3476 489972 3528
rect 490564 3476 490616 3528
rect 505376 3476 505428 3528
rect 507124 3476 507176 3528
rect 523040 3476 523092 3528
rect 523684 3476 523736 3528
rect 526720 3476 526772 3528
rect 526996 3476 527048 3528
rect 544384 3476 544436 3528
rect 544660 3476 544712 3528
rect 563244 3476 563296 3528
rect 563428 3476 563480 3528
rect 583392 3476 583444 3528
rect 479340 3408 479392 3460
rect 438676 3340 438728 3392
rect 449808 3340 449860 3392
rect 455236 3340 455288 3392
rect 467472 3340 467524 3392
rect 469588 3340 469640 3392
rect 447508 3272 447560 3324
rect 459192 3272 459244 3324
rect 52552 3204 52604 3256
rect 67732 3204 67784 3256
rect 72608 3204 72660 3256
rect 86500 3204 86552 3256
rect 90364 3204 90416 3256
rect 103060 3204 103112 3256
rect 106924 3204 106976 3256
rect 118516 3204 118568 3256
rect 181444 3204 181496 3256
rect 188068 3204 188120 3256
rect 201500 3204 201552 3256
rect 206836 3204 206888 3256
rect 210976 3204 211028 3256
rect 215668 3204 215720 3256
rect 331588 3204 331640 3256
rect 335084 3204 335136 3256
rect 356980 3204 357032 3256
rect 362316 3204 362368 3256
rect 440884 3204 440936 3256
rect 452108 3204 452160 3256
rect 454132 3204 454184 3256
rect 466276 3204 466328 3256
rect 24216 3136 24268 3188
rect 41236 3136 41288 3188
rect 47860 3136 47912 3188
rect 63316 3136 63368 3188
rect 65524 3136 65576 3188
rect 79876 3136 79928 3188
rect 85672 3136 85724 3188
rect 98276 3136 98328 3188
rect 182548 3136 182600 3188
rect 189172 3136 189224 3188
rect 192024 3136 192076 3188
rect 198004 3136 198056 3188
rect 203892 3136 203944 3188
rect 209044 3136 209096 3188
rect 213368 3136 213420 3188
rect 217876 3136 217928 3188
rect 223948 3136 224000 3188
rect 227812 3136 227864 3188
rect 229836 3136 229888 3188
rect 233332 3136 233384 3188
rect 246396 3136 246448 3188
rect 248788 3136 248840 3188
rect 298468 3136 298520 3188
rect 299664 3136 299716 3188
rect 322756 3136 322808 3188
rect 325608 3136 325660 3188
rect 341524 3136 341576 3188
rect 345756 3136 345808 3188
rect 348148 3136 348200 3188
rect 352840 3136 352892 3188
rect 360292 3136 360344 3188
rect 365812 3136 365864 3188
rect 370228 3136 370280 3188
rect 376484 3136 376536 3188
rect 376852 3136 376904 3188
rect 383568 3136 383620 3188
rect 384580 3136 384632 3188
rect 391848 3136 391900 3188
rect 393412 3136 393464 3188
rect 401324 3136 401376 3188
rect 449716 3136 449768 3188
rect 461584 3136 461636 3188
rect 472900 3272 472952 3324
rect 486424 3408 486476 3460
rect 489460 3408 489512 3460
rect 504180 3408 504232 3460
rect 506020 3408 506072 3460
rect 521844 3408 521896 3460
rect 522580 3408 522632 3460
rect 539600 3408 539652 3460
rect 542452 3408 542504 3460
rect 560852 3408 560904 3460
rect 561220 3408 561272 3460
rect 581000 3408 581052 3460
rect 482836 3340 482888 3392
rect 486148 3340 486200 3392
rect 500592 3340 500644 3392
rect 500776 3340 500828 3392
rect 515956 3340 516008 3392
rect 516048 3340 516100 3392
rect 532516 3340 532568 3392
rect 532608 3340 532660 3392
rect 550272 3340 550324 3392
rect 554596 3340 554648 3392
rect 573916 3340 573968 3392
rect 19432 3068 19484 3120
rect 36820 3068 36872 3120
rect 44272 3068 44324 3120
rect 60004 3068 60056 3120
rect 60832 3068 60884 3120
rect 75460 3068 75512 3120
rect 102232 3068 102284 3120
rect 114100 3068 114152 3120
rect 164884 3068 164936 3120
rect 172612 3068 172664 3120
rect 184940 3068 184992 3120
rect 191380 3068 191432 3120
rect 195612 3068 195664 3120
rect 201316 3068 201368 3120
rect 205088 3068 205140 3120
rect 210148 3068 210200 3120
rect 215668 3068 215720 3120
rect 220084 3068 220136 3120
rect 221556 3068 221608 3120
rect 225604 3068 225656 3120
rect 226340 3068 226392 3120
rect 230020 3068 230072 3120
rect 231032 3068 231084 3120
rect 234436 3068 234488 3120
rect 234620 3068 234672 3120
rect 237748 3068 237800 3120
rect 238116 3068 238168 3120
rect 241060 3068 241112 3120
rect 241704 3068 241756 3120
rect 244372 3068 244424 3120
rect 247592 3068 247644 3120
rect 249892 3068 249944 3120
rect 249984 3068 250036 3120
rect 252100 3068 252152 3120
rect 252376 3068 252428 3120
rect 254308 3068 254360 3120
rect 254676 3068 254728 3120
rect 256516 3068 256568 3120
rect 257068 3068 257120 3120
rect 258724 3068 258776 3120
rect 259460 3068 259512 3120
rect 260932 3068 260984 3120
rect 261760 3068 261812 3120
rect 263140 3068 263192 3120
rect 264152 3068 264204 3120
rect 265348 3068 265400 3120
rect 271236 3068 271288 3120
rect 271972 3068 272024 3120
rect 300676 3068 300728 3120
rect 301964 3068 302016 3120
rect 302884 3068 302936 3120
rect 304356 3068 304408 3120
rect 305092 3068 305144 3120
rect 306748 3068 306800 3120
rect 307300 3068 307352 3120
rect 309048 3068 309100 3120
rect 311716 3068 311768 3120
rect 313832 3068 313884 3120
rect 315028 3068 315080 3120
rect 317328 3068 317380 3120
rect 319444 3068 319496 3120
rect 322112 3068 322164 3120
rect 324964 3068 325016 3120
rect 328000 3068 328052 3120
rect 328276 3068 328328 3120
rect 331588 3068 331640 3120
rect 332692 3068 332744 3120
rect 336280 3068 336332 3120
rect 337108 3068 337160 3120
rect 340972 3068 341024 3120
rect 345940 3068 345992 3120
rect 350448 3068 350500 3120
rect 359188 3068 359240 3120
rect 364616 3068 364668 3120
rect 369124 3068 369176 3120
rect 375288 3068 375340 3120
rect 379060 3068 379112 3120
rect 385960 3068 386012 3120
rect 386788 3068 386840 3120
rect 394240 3068 394292 3120
rect 403348 3068 403400 3120
rect 411904 3068 411956 3120
rect 470692 3068 470744 3120
rect 484032 3272 484084 3324
rect 487252 3272 487304 3324
rect 501788 3272 501840 3324
rect 501880 3272 501932 3324
rect 517152 3272 517204 3324
rect 524788 3272 524840 3324
rect 492772 3204 492824 3256
rect 507676 3204 507728 3256
rect 509332 3204 509384 3256
rect 525432 3204 525484 3256
rect 526720 3272 526772 3324
rect 540796 3272 540848 3324
rect 541992 3204 542044 3256
rect 485044 3136 485096 3188
rect 499396 3136 499448 3188
rect 517060 3136 517112 3188
rect 533712 3136 533764 3188
rect 540244 3136 540296 3188
rect 558552 3272 558604 3324
rect 546868 3204 546920 3256
rect 565636 3204 565688 3256
rect 480628 3068 480680 3120
rect 494704 3068 494756 3120
rect 503812 3068 503864 3120
rect 519544 3068 519596 3120
rect 531412 3068 531464 3120
rect 549076 3068 549128 3120
rect 18236 3000 18288 3052
rect 35716 3000 35768 3052
rect 69112 3000 69164 3052
rect 83188 3000 83240 3052
rect 142436 3000 142488 3052
rect 151636 3000 151688 3052
rect 151820 3000 151872 3052
rect 160468 3000 160520 3052
rect 166080 3000 166132 3052
rect 173716 3000 173768 3052
rect 186136 3000 186188 3052
rect 192484 3000 192536 3052
rect 196808 3000 196860 3052
rect 202420 3000 202472 3052
rect 207388 3000 207440 3052
rect 212356 3000 212408 3052
rect 216864 3000 216916 3052
rect 221188 3000 221240 3052
rect 222752 3000 222804 3052
rect 226708 3000 226760 3052
rect 227536 3000 227588 3052
rect 231124 3000 231176 3052
rect 233424 3000 233476 3052
rect 236644 3000 236696 3052
rect 237012 3000 237064 3052
rect 239956 3000 240008 3052
rect 240508 3000 240560 3052
rect 243268 3000 243320 3052
rect 244096 3000 244148 3052
rect 246580 3000 246632 3052
rect 248788 3000 248840 3052
rect 250996 3000 251048 3052
rect 251180 3000 251232 3052
rect 253204 3000 253256 3052
rect 253480 3000 253532 3052
rect 255412 3000 255464 3052
rect 255872 3000 255924 3052
rect 257620 3000 257672 3052
rect 258264 3000 258316 3052
rect 259828 3000 259880 3052
rect 260656 3000 260708 3052
rect 262036 3000 262088 3052
rect 262956 3000 263008 3052
rect 264244 3000 264296 3052
rect 267740 3000 267792 3052
rect 268660 3000 268712 3052
rect 291844 3000 291896 3052
rect 292580 3000 292632 3052
rect 294052 3000 294104 3052
rect 294880 3000 294932 3052
rect 295156 3000 295208 3052
rect 296076 3000 296128 3052
rect 296260 3000 296312 3052
rect 297272 3000 297324 3052
rect 297364 3000 297416 3052
rect 298468 3000 298520 3052
rect 299572 3000 299624 3052
rect 300768 3000 300820 3052
rect 301780 3000 301832 3052
rect 303160 3000 303212 3052
rect 303988 3000 304040 3052
rect 305552 3000 305604 3052
rect 306196 3000 306248 3052
rect 307944 3000 307996 3052
rect 308404 3000 308456 3052
rect 310244 3000 310296 3052
rect 310612 3000 310664 3052
rect 312636 3000 312688 3052
rect 313924 3000 313976 3052
rect 316224 3000 316276 3052
rect 317236 3000 317288 3052
rect 319720 3000 319772 3052
rect 320548 3000 320600 3052
rect 323308 3000 323360 3052
rect 326068 3000 326120 3052
rect 329196 3000 329248 3052
rect 330484 3000 330536 3052
rect 333888 3000 333940 3052
rect 336004 3000 336056 3052
rect 339868 3000 339920 3052
rect 340420 3000 340472 3052
rect 344560 3000 344612 3052
rect 347044 3000 347096 3052
rect 351644 3000 351696 3052
rect 354772 3000 354824 3052
rect 359924 3000 359976 3052
rect 364708 3000 364760 3052
rect 370596 3000 370648 3052
rect 374644 3000 374696 3052
rect 381176 3000 381228 3052
rect 387892 3000 387944 3052
rect 395344 3000 395396 3052
rect 396724 3000 396776 3052
rect 404820 3000 404872 3052
rect 508228 3000 508280 3052
rect 524236 3000 524288 3052
rect 541348 3000 541400 3052
rect 559748 3136 559800 3188
rect 25320 2932 25372 2984
rect 42340 2932 42392 2984
rect 59636 2932 59688 2984
rect 74356 2932 74408 2984
rect 162492 2932 162544 2984
rect 170404 2932 170456 2984
rect 171968 2932 172020 2984
rect 179236 2932 179288 2984
rect 183744 2932 183796 2984
rect 190276 2932 190328 2984
rect 194416 2932 194468 2984
rect 200212 2932 200264 2984
rect 200304 2932 200356 2984
rect 205732 2932 205784 2984
rect 206192 2932 206244 2984
rect 211252 2932 211304 2984
rect 214472 2932 214524 2984
rect 218980 2932 219032 2984
rect 220452 2932 220504 2984
rect 224500 2932 224552 2984
rect 225144 2932 225196 2984
rect 228916 2932 228968 2984
rect 232228 2932 232280 2984
rect 235540 2932 235592 2984
rect 239312 2932 239364 2984
rect 242164 2932 242216 2984
rect 245200 2932 245252 2984
rect 247684 2932 247736 2984
rect 316132 2932 316184 2984
rect 318524 2932 318576 2984
rect 323860 2932 323912 2984
rect 326804 2932 326856 2984
rect 327172 2932 327224 2984
rect 330392 2932 330444 2984
rect 333796 2932 333848 2984
rect 337476 2932 337528 2984
rect 338212 2932 338264 2984
rect 342168 2932 342220 2984
rect 342628 2932 342680 2984
rect 346952 2932 347004 2984
rect 351460 2932 351512 2984
rect 356336 2932 356388 2984
rect 361396 2932 361448 2984
rect 367008 2932 367060 2984
rect 368020 2932 368072 2984
rect 374092 2932 374144 2984
rect 377956 2932 378008 2984
rect 384764 2932 384816 2984
rect 385684 2932 385736 2984
rect 393044 2932 393096 2984
rect 394516 2932 394568 2984
rect 402520 2932 402572 2984
rect 547972 2932 548024 2984
rect 566832 3068 566884 3120
rect 27712 2864 27764 2916
rect 44548 2864 44600 2916
rect 155408 2864 155460 2916
rect 163780 2864 163832 2916
rect 173164 2864 173216 2916
rect 180340 2864 180392 2916
rect 190828 2864 190880 2916
rect 196900 2864 196952 2916
rect 202696 2864 202748 2916
rect 207940 2864 207992 2916
rect 212172 2864 212224 2916
rect 216772 2864 216824 2916
rect 235816 2864 235868 2916
rect 238852 2864 238904 2916
rect 242900 2864 242952 2916
rect 245476 2864 245528 2916
rect 265348 2864 265400 2916
rect 266452 2864 266504 2916
rect 268844 2864 268896 2916
rect 269764 2864 269816 2916
rect 329380 2864 329432 2916
rect 332692 2864 332744 2916
rect 339316 2864 339368 2916
rect 343364 2864 343416 2916
rect 350356 2864 350408 2916
rect 355232 2864 355284 2916
rect 355876 2864 355928 2916
rect 361120 2864 361172 2916
rect 375748 2864 375800 2916
rect 382372 2864 382424 2916
rect 35992 2796 36044 2848
rect 52276 2796 52328 2848
rect 209780 2796 209832 2848
rect 214564 2796 214616 2848
rect 309508 2796 309560 2848
rect 311440 2796 311492 2848
rect 312820 2796 312872 2848
rect 315028 2796 315080 2848
rect 318340 2796 318392 2848
rect 320916 2796 320968 2848
rect 321652 2796 321704 2848
rect 324412 2796 324464 2848
rect 358084 2796 358136 2848
rect 363512 2796 363564 2848
rect 366916 2796 366968 2848
rect 372896 2796 372948 2848
rect 474740 2796 474792 2848
rect 475752 2796 475804 2848
rect 525800 2796 525852 2848
rect 526628 2796 526680 2848
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218072 703582 218836 703610
rect 8128 700330 8156 703520
rect 8116 700324 8168 700330
rect 8116 700266 8168 700272
rect 13912 700324 13964 700330
rect 13912 700266 13964 700272
rect 3422 697368 3478 697377
rect 3422 697303 3478 697312
rect 3436 684457 3464 697303
rect 13924 692594 13952 700266
rect 24320 699718 24348 703520
rect 40512 700398 40540 703520
rect 56796 700534 56824 703520
rect 56784 700528 56836 700534
rect 56784 700470 56836 700476
rect 61384 700528 61436 700534
rect 61384 700470 61436 700476
rect 40500 700392 40552 700398
rect 40500 700334 40552 700340
rect 44180 700392 44232 700398
rect 44180 700334 44232 700340
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 28264 699712 28316 699718
rect 28264 699654 28316 699660
rect 28276 695502 28304 699654
rect 28264 695496 28316 695502
rect 28264 695438 28316 695444
rect 30196 695496 30248 695502
rect 30196 695438 30248 695444
rect 13924 692566 14398 692594
rect 30208 692580 30236 695438
rect 44192 694210 44220 700334
rect 44180 694204 44232 694210
rect 44180 694146 44232 694152
rect 46020 694204 46072 694210
rect 46020 694146 46072 694152
rect 46032 692580 46060 694146
rect 61396 692594 61424 700470
rect 72988 699718 73016 703520
rect 89180 700738 89208 703520
rect 105464 700942 105492 703520
rect 105452 700936 105504 700942
rect 105452 700878 105504 700884
rect 109040 700936 109092 700942
rect 109040 700878 109092 700884
rect 89168 700732 89220 700738
rect 89168 700674 89220 700680
rect 93032 700732 93084 700738
rect 93032 700674 93084 700680
rect 72976 699712 73028 699718
rect 72976 699654 73028 699660
rect 76104 699712 76156 699718
rect 76104 699654 76156 699660
rect 76116 695502 76144 699654
rect 76104 695496 76156 695502
rect 76104 695438 76156 695444
rect 77668 695496 77720 695502
rect 77668 695438 77720 695444
rect 61396 692566 61870 692594
rect 77680 692580 77708 695438
rect 93044 692594 93072 700674
rect 109052 692594 109080 700878
rect 121656 694210 121684 703520
rect 137848 699718 137876 703520
rect 154132 702434 154160 703520
rect 170324 702434 170352 703520
rect 153212 702406 154160 702434
rect 169772 702406 170352 702434
rect 137836 699712 137888 699718
rect 137836 699654 137888 699660
rect 140780 699712 140832 699718
rect 140780 699654 140832 699660
rect 121644 694204 121696 694210
rect 121644 694146 121696 694152
rect 125140 694204 125192 694210
rect 125140 694146 125192 694152
rect 93044 692566 93518 692594
rect 109052 692566 109342 692594
rect 125152 692580 125180 694146
rect 140792 692594 140820 699654
rect 153212 695502 153240 702406
rect 153200 695496 153252 695502
rect 153200 695438 153252 695444
rect 156788 695496 156840 695502
rect 156788 695438 156840 695444
rect 140792 692566 140990 692594
rect 156800 692580 156828 695438
rect 169772 694210 169800 702406
rect 186516 695502 186544 703520
rect 202800 703050 202828 703520
rect 201500 703044 201552 703050
rect 201500 702986 201552 702992
rect 202788 703044 202840 703050
rect 202788 702986 202840 702992
rect 201512 695502 201540 702986
rect 186504 695496 186556 695502
rect 186504 695438 186556 695444
rect 188436 695496 188488 695502
rect 188436 695438 188488 695444
rect 201500 695496 201552 695502
rect 201500 695438 201552 695444
rect 204260 695496 204312 695502
rect 204260 695438 204312 695444
rect 169760 694204 169812 694210
rect 169760 694146 169812 694152
rect 172612 694204 172664 694210
rect 172612 694146 172664 694152
rect 172624 692580 172652 694146
rect 188448 692580 188476 695438
rect 204272 692580 204300 695438
rect 218072 694210 218100 703582
rect 218808 703474 218836 703582
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 218992 703474 219020 703520
rect 218808 703446 219020 703474
rect 235184 702434 235212 703520
rect 251468 702434 251496 703520
rect 235184 702406 235488 702434
rect 218060 694204 218112 694210
rect 218060 694146 218112 694152
rect 220084 694204 220136 694210
rect 220084 694146 220136 694152
rect 220096 692580 220124 694146
rect 235460 692594 235488 702406
rect 251284 702406 251496 702434
rect 251284 692594 251312 702406
rect 267660 692594 267688 703520
rect 283852 702434 283880 703520
rect 235460 692566 235934 692594
rect 251284 692566 251758 692594
rect 267582 692566 267688 692594
rect 282932 702406 283880 702434
rect 282932 692594 282960 702406
rect 300136 699718 300164 703520
rect 316328 699718 316356 703520
rect 332520 699718 332548 703520
rect 348804 699718 348832 703520
rect 364996 699718 365024 703520
rect 381188 699718 381216 703520
rect 397472 699718 397500 703520
rect 413664 699718 413692 703520
rect 429856 699718 429884 703520
rect 446140 699718 446168 703520
rect 298744 699712 298796 699718
rect 298744 699654 298796 699660
rect 300124 699712 300176 699718
rect 300124 699654 300176 699660
rect 314660 699712 314712 699718
rect 314660 699654 314712 699660
rect 316316 699712 316368 699718
rect 316316 699654 316368 699660
rect 330392 699712 330444 699718
rect 330392 699654 330444 699660
rect 332508 699712 332560 699718
rect 332508 699654 332560 699660
rect 346400 699712 346452 699718
rect 346400 699654 346452 699660
rect 348792 699712 348844 699718
rect 348792 699654 348844 699660
rect 362040 699712 362092 699718
rect 362040 699654 362092 699660
rect 364984 699712 365036 699718
rect 364984 699654 365036 699660
rect 378140 699712 378192 699718
rect 378140 699654 378192 699660
rect 381176 699712 381228 699718
rect 381176 699654 381228 699660
rect 393688 699712 393740 699718
rect 393688 699654 393740 699660
rect 397460 699712 397512 699718
rect 397460 699654 397512 699660
rect 409880 699712 409932 699718
rect 409880 699654 409932 699660
rect 413652 699712 413704 699718
rect 413652 699654 413704 699660
rect 425336 699712 425388 699718
rect 425336 699654 425388 699660
rect 429844 699712 429896 699718
rect 429844 699654 429896 699660
rect 441620 699712 441672 699718
rect 441620 699654 441672 699660
rect 446128 699712 446180 699718
rect 446128 699654 446180 699660
rect 298756 692594 298784 699654
rect 314672 692594 314700 699654
rect 330404 692594 330432 699654
rect 346412 692594 346440 699654
rect 362052 692594 362080 699654
rect 378152 692594 378180 699654
rect 393700 692594 393728 699654
rect 409892 692594 409920 699654
rect 425348 692594 425376 699654
rect 282932 692566 283406 692594
rect 298756 692566 299230 692594
rect 314672 692566 315054 692594
rect 330404 692566 330878 692594
rect 346412 692566 346702 692594
rect 362052 692566 362526 692594
rect 378152 692566 378350 692594
rect 393700 692566 394174 692594
rect 409892 692566 409998 692594
rect 425348 692566 425822 692594
rect 441632 692580 441660 699654
rect 462332 694210 462360 703520
rect 478524 702434 478552 703520
rect 477512 702406 478552 702434
rect 477512 695434 477540 702406
rect 473268 695428 473320 695434
rect 473268 695370 473320 695376
rect 477500 695428 477552 695434
rect 477500 695370 477552 695376
rect 457444 694204 457496 694210
rect 457444 694146 457496 694152
rect 462320 694204 462372 694210
rect 462320 694146 462372 694152
rect 457456 692580 457484 694146
rect 473280 692580 473308 695370
rect 494072 694822 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510632 703582 510844 703610
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 489092 694816 489144 694822
rect 489092 694758 489144 694764
rect 494060 694816 494112 694822
rect 494060 694758 494112 694764
rect 489104 692580 489132 694758
rect 510632 694210 510660 703582
rect 510816 703474 510844 703582
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 511000 703474 511028 703520
rect 510816 703446 511028 703474
rect 527192 695502 527220 703520
rect 543476 702434 543504 703520
rect 559668 702434 559696 703520
rect 542372 702406 543504 702434
rect 558932 702406 559696 702434
rect 520740 695496 520792 695502
rect 520740 695438 520792 695444
rect 527180 695496 527232 695502
rect 527180 695438 527232 695444
rect 504916 694204 504968 694210
rect 504916 694146 504968 694152
rect 510620 694204 510672 694210
rect 510620 694146 510672 694152
rect 504928 692580 504956 694146
rect 520752 692580 520780 695438
rect 542372 694822 542400 702406
rect 536564 694816 536616 694822
rect 536564 694758 536616 694764
rect 542360 694816 542412 694822
rect 542360 694758 542412 694764
rect 536576 692580 536604 694758
rect 558932 694210 558960 702406
rect 575860 699718 575888 703520
rect 574100 699712 574152 699718
rect 574100 699654 574152 699660
rect 575848 699712 575900 699718
rect 575848 699654 575900 699660
rect 574112 695298 574140 699654
rect 578882 697232 578938 697241
rect 578882 697167 578938 697176
rect 568212 695292 568264 695298
rect 568212 695234 568264 695240
rect 574100 695292 574152 695298
rect 574100 695234 574152 695240
rect 552388 694204 552440 694210
rect 552388 694146 552440 694152
rect 558920 694204 558972 694210
rect 558920 694146 558972 694152
rect 552400 692580 552428 694146
rect 568224 692580 568252 695234
rect 578896 685273 578924 697167
rect 578882 685264 578938 685273
rect 578882 685199 578938 685208
rect 3422 684448 3478 684457
rect 3422 684383 3478 684392
rect 3606 684312 3662 684321
rect 3606 684247 3662 684256
rect 3620 671809 3648 684247
rect 580262 683904 580318 683913
rect 580262 683839 580318 683848
rect 580276 672994 580304 683839
rect 578332 672988 578384 672994
rect 578332 672930 578384 672936
rect 580264 672988 580316 672994
rect 580264 672930 580316 672936
rect 578344 672353 578372 672930
rect 578330 672344 578386 672353
rect 578330 672279 578386 672288
rect 3606 671800 3662 671809
rect 3606 671735 3662 671744
rect 3422 671256 3478 671265
rect 3422 671191 3478 671200
rect 3436 659161 3464 671191
rect 580262 670712 580318 670721
rect 580262 670647 580318 670656
rect 580276 659462 580304 670647
rect 578516 659456 578568 659462
rect 578514 659424 578516 659433
rect 580264 659456 580316 659462
rect 578568 659424 578570 659433
rect 580264 659398 580316 659404
rect 578514 659359 578570 659368
rect 3422 659152 3478 659161
rect 3422 659087 3478 659096
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 646513 3464 658135
rect 580262 657384 580318 657393
rect 580262 657319 580318 657328
rect 580276 647018 580304 657319
rect 578332 647012 578384 647018
rect 578332 646954 578384 646960
rect 580264 647012 580316 647018
rect 580264 646954 580316 646960
rect 578344 646513 578372 646954
rect 3422 646504 3478 646513
rect 3422 646439 3478 646448
rect 578330 646504 578386 646513
rect 578330 646439 578386 646448
rect 3422 645144 3478 645153
rect 3422 645079 3478 645088
rect 3436 633865 3464 645079
rect 578882 644056 578938 644065
rect 578882 643991 578938 644000
rect 3422 633856 3478 633865
rect 3422 633791 3478 633800
rect 578896 633593 578924 643991
rect 578882 633584 578938 633593
rect 578882 633519 578938 633528
rect 3422 632088 3478 632097
rect 3422 632023 3478 632032
rect 3436 621217 3464 632023
rect 580262 630864 580318 630873
rect 580262 630799 580318 630808
rect 3422 621208 3478 621217
rect 3422 621143 3478 621152
rect 580276 620974 580304 630799
rect 578332 620968 578384 620974
rect 578332 620910 578384 620916
rect 580264 620968 580316 620974
rect 580264 620910 580316 620916
rect 578344 620673 578372 620910
rect 578330 620664 578386 620673
rect 578330 620599 578386 620608
rect 3422 619168 3478 619177
rect 3422 619103 3478 619112
rect 3436 608569 3464 619103
rect 578882 617536 578938 617545
rect 578882 617471 578938 617480
rect 3422 608560 3478 608569
rect 3422 608495 3478 608504
rect 578896 607753 578924 617471
rect 578882 607744 578938 607753
rect 578882 607679 578938 607688
rect 3422 606112 3478 606121
rect 3422 606047 3478 606056
rect 3436 595921 3464 606047
rect 578882 604208 578938 604217
rect 578882 604143 578938 604152
rect 3422 595912 3478 595921
rect 3422 595847 3478 595856
rect 578896 594833 578924 604143
rect 578882 594824 578938 594833
rect 578882 594759 578938 594768
rect 3422 593056 3478 593065
rect 3422 592991 3478 593000
rect 3436 583273 3464 592991
rect 578882 591016 578938 591025
rect 578882 590951 578938 590960
rect 3422 583264 3478 583273
rect 3422 583199 3478 583208
rect 578896 581913 578924 590951
rect 578882 581904 578938 581913
rect 578882 581839 578938 581848
rect 3422 580000 3478 580009
rect 3422 579935 3478 579944
rect 3436 570625 3464 579935
rect 578882 577688 578938 577697
rect 578882 577623 578938 577632
rect 3422 570616 3478 570625
rect 3422 570551 3478 570560
rect 578896 568993 578924 577623
rect 578882 568984 578938 568993
rect 578882 568919 578938 568928
rect 3054 566944 3110 566953
rect 3054 566879 3110 566888
rect 3068 557977 3096 566879
rect 578882 564360 578938 564369
rect 578882 564295 578938 564304
rect 3054 557968 3110 557977
rect 3054 557903 3110 557912
rect 578896 556073 578924 564295
rect 578882 556064 578938 556073
rect 578882 555999 578938 556008
rect 3422 553888 3478 553897
rect 3422 553823 3478 553832
rect 3436 545329 3464 553823
rect 578882 551168 578938 551177
rect 578882 551103 578938 551112
rect 3422 545320 3478 545329
rect 3422 545255 3478 545264
rect 578896 543153 578924 551103
rect 578882 543144 578938 543153
rect 578882 543079 578938 543088
rect 2962 540832 3018 540841
rect 2962 540767 3018 540776
rect 2976 532681 3004 540767
rect 579526 537840 579582 537849
rect 579526 537775 579582 537784
rect 2962 532672 3018 532681
rect 2962 532607 3018 532616
rect 579540 530233 579568 537775
rect 579526 530224 579582 530233
rect 579526 530159 579582 530168
rect 2962 527912 3018 527921
rect 2962 527847 3018 527856
rect 2976 520033 3004 527847
rect 578882 524512 578938 524521
rect 578882 524447 578938 524456
rect 2962 520024 3018 520033
rect 2962 519959 3018 519968
rect 578896 517313 578924 524447
rect 578882 517304 578938 517313
rect 578882 517239 578938 517248
rect 3422 514856 3478 514865
rect 3422 514791 3478 514800
rect 3436 507385 3464 514791
rect 580538 511320 580594 511329
rect 580538 511255 580594 511264
rect 580552 510678 580580 511255
rect 578240 510672 578292 510678
rect 578240 510614 578292 510620
rect 580540 510672 580592 510678
rect 580540 510614 580592 510620
rect 3422 507376 3478 507385
rect 3422 507311 3478 507320
rect 578252 504393 578280 510614
rect 578238 504384 578294 504393
rect 578238 504319 578294 504328
rect 3054 501800 3110 501809
rect 3054 501735 3110 501744
rect 3068 494737 3096 501735
rect 579526 497992 579582 498001
rect 579526 497927 579582 497936
rect 3054 494728 3110 494737
rect 3054 494663 3110 494672
rect 579540 491473 579568 497927
rect 579526 491464 579582 491473
rect 579526 491399 579582 491408
rect 2962 488744 3018 488753
rect 2962 488679 3018 488688
rect 2976 482089 3004 488679
rect 578882 484664 578938 484673
rect 578882 484599 578938 484608
rect 2962 482080 3018 482089
rect 2962 482015 3018 482024
rect 578896 478553 578924 484599
rect 578882 478544 578938 478553
rect 578882 478479 578938 478488
rect 3422 475688 3478 475697
rect 3422 475623 3478 475632
rect 3436 469441 3464 475623
rect 579802 471472 579858 471481
rect 579802 471407 579858 471416
rect 579816 471034 579844 471407
rect 578240 471028 578292 471034
rect 578240 470970 578292 470976
rect 579804 471028 579856 471034
rect 579804 470970 579856 470976
rect 3422 469432 3478 469441
rect 3422 469367 3478 469376
rect 578252 465633 578280 470970
rect 578238 465624 578294 465633
rect 578238 465559 578294 465568
rect 2962 462632 3018 462641
rect 2962 462567 3018 462576
rect 2976 456793 3004 462567
rect 579526 458144 579582 458153
rect 579526 458079 579582 458088
rect 2962 456784 3018 456793
rect 2962 456719 3018 456728
rect 579540 452713 579568 458079
rect 579526 452704 579582 452713
rect 579526 452639 579582 452648
rect 3054 449576 3110 449585
rect 3054 449511 3110 449520
rect 3068 444145 3096 449511
rect 578882 444816 578938 444825
rect 578882 444751 578938 444760
rect 3054 444136 3110 444145
rect 3054 444071 3110 444080
rect 578896 439793 578924 444751
rect 578882 439784 578938 439793
rect 578882 439719 578938 439728
rect 3422 436656 3478 436665
rect 3422 436591 3478 436600
rect 3436 431497 3464 436591
rect 579526 431624 579582 431633
rect 579526 431559 579582 431568
rect 3422 431488 3478 431497
rect 3422 431423 3478 431432
rect 579540 426873 579568 431559
rect 579526 426864 579582 426873
rect 579526 426799 579582 426808
rect 2962 423600 3018 423609
rect 2962 423535 3018 423544
rect 2976 418849 3004 423535
rect 2962 418840 3018 418849
rect 2962 418775 3018 418784
rect 579526 418296 579582 418305
rect 579526 418231 579582 418240
rect 579540 413953 579568 418231
rect 579526 413944 579582 413953
rect 579526 413879 579582 413888
rect 3054 410544 3110 410553
rect 3054 410479 3110 410488
rect 3068 406201 3096 410479
rect 3054 406192 3110 406201
rect 3054 406127 3110 406136
rect 580354 404968 580410 404977
rect 580354 404903 580410 404912
rect 580368 404394 580396 404903
rect 578240 404388 578292 404394
rect 578240 404330 578292 404336
rect 580356 404388 580408 404394
rect 580356 404330 580408 404336
rect 578252 401033 578280 404330
rect 578238 401024 578294 401033
rect 578238 400959 578294 400968
rect 2778 397488 2834 397497
rect 2778 397423 2834 397432
rect 2792 393553 2820 397423
rect 2778 393544 2834 393553
rect 2778 393479 2834 393488
rect 579618 391776 579674 391785
rect 579618 391711 579674 391720
rect 579526 388104 579582 388113
rect 579632 388090 579660 391711
rect 579582 388062 579660 388090
rect 579526 388039 579582 388048
rect 3054 384432 3110 384441
rect 3054 384367 3110 384376
rect 3068 380905 3096 384367
rect 3054 380896 3110 380905
rect 3054 380831 3110 380840
rect 579526 378448 579582 378457
rect 579526 378383 579582 378392
rect 579540 375193 579568 378383
rect 579526 375184 579582 375193
rect 579526 375119 579582 375128
rect 3054 371376 3110 371385
rect 3054 371311 3110 371320
rect 3068 368257 3096 371311
rect 3054 368248 3110 368257
rect 3054 368183 3110 368192
rect 580906 365120 580962 365129
rect 580906 365055 580962 365064
rect 580920 362778 580948 365055
rect 578332 362772 578384 362778
rect 578332 362714 578384 362720
rect 580908 362772 580960 362778
rect 580908 362714 580960 362720
rect 578344 362273 578372 362714
rect 578330 362264 578386 362273
rect 578330 362199 578386 362208
rect 3054 358456 3110 358465
rect 3054 358391 3110 358400
rect 3068 355609 3096 358391
rect 3054 355600 3110 355609
rect 3054 355535 3110 355544
rect 579618 351928 579674 351937
rect 579618 351863 579674 351872
rect 579526 349344 579582 349353
rect 579632 349330 579660 351863
rect 579582 349302 579660 349330
rect 579526 349279 579582 349288
rect 3054 345400 3110 345409
rect 3054 345335 3110 345344
rect 3068 342961 3096 345335
rect 3054 342952 3110 342961
rect 3054 342887 3110 342896
rect 579618 338600 579674 338609
rect 579618 338535 579674 338544
rect 579526 336424 579582 336433
rect 579632 336410 579660 338535
rect 579582 336382 579660 336410
rect 579526 336359 579582 336368
rect 3054 332344 3110 332353
rect 3054 332279 3110 332288
rect 3068 330313 3096 332279
rect 3054 330304 3110 330313
rect 3054 330239 3110 330248
rect 579618 325272 579674 325281
rect 579618 325207 579674 325216
rect 579526 323504 579582 323513
rect 579632 323490 579660 325207
rect 579582 323462 579660 323490
rect 579526 323439 579582 323448
rect 3054 319288 3110 319297
rect 3054 319223 3110 319232
rect 3068 317665 3096 319223
rect 3054 317656 3110 317665
rect 3054 317591 3110 317600
rect 579618 312080 579674 312089
rect 579618 312015 579674 312024
rect 579526 310584 579582 310593
rect 579632 310570 579660 312015
rect 579582 310542 579660 310570
rect 579526 310519 579582 310528
rect 3054 306232 3110 306241
rect 3054 306167 3110 306176
rect 3068 305017 3096 306167
rect 3054 305008 3110 305017
rect 3054 304943 3110 304952
rect 579618 298752 579674 298761
rect 579618 298687 579674 298696
rect 579526 297664 579582 297673
rect 579632 297650 579660 298687
rect 579582 297622 579660 297650
rect 579526 297599 579582 297608
rect 3054 293176 3110 293185
rect 3054 293111 3110 293120
rect 3068 292369 3096 293111
rect 3054 292360 3110 292369
rect 3054 292295 3110 292304
rect 3054 229120 3110 229129
rect 3054 229055 3110 229064
rect 3068 228041 3096 229055
rect 3054 228032 3110 228041
rect 3054 227967 3110 227976
rect 578514 220144 578570 220153
rect 578514 220079 578570 220088
rect 578528 219774 578556 220079
rect 578516 219768 578568 219774
rect 578516 219710 578568 219716
rect 580908 219768 580960 219774
rect 580908 219710 580960 219716
rect 580920 219065 580948 219710
rect 580906 219056 580962 219065
rect 580906 218991 580962 219000
rect 3054 216472 3110 216481
rect 3054 216407 3110 216416
rect 3068 214985 3096 216407
rect 3054 214976 3110 214985
rect 3054 214911 3110 214920
rect 579526 207224 579582 207233
rect 579582 207182 579660 207210
rect 579526 207159 579582 207168
rect 579632 205737 579660 207182
rect 579618 205728 579674 205737
rect 579618 205663 579674 205672
rect 3054 203824 3110 203833
rect 3054 203759 3110 203768
rect 3068 201929 3096 203759
rect 3054 201920 3110 201929
rect 3054 201855 3110 201864
rect 579526 194304 579582 194313
rect 579582 194262 579660 194290
rect 579526 194239 579582 194248
rect 579632 192545 579660 194262
rect 579618 192536 579674 192545
rect 579618 192471 579674 192480
rect 2962 191176 3018 191185
rect 2962 191111 3018 191120
rect 2976 188873 3004 191111
rect 2962 188864 3018 188873
rect 2962 188799 3018 188808
rect 578330 181384 578386 181393
rect 578330 181319 578332 181328
rect 578384 181319 578386 181328
rect 580540 181348 580592 181354
rect 578332 181290 578384 181296
rect 580540 181290 580592 181296
rect 580552 179217 580580 181290
rect 580538 179208 580594 179217
rect 580538 179143 580594 179152
rect 2962 178528 3018 178537
rect 2962 178463 3018 178472
rect 2976 175953 3004 178463
rect 2962 175944 3018 175953
rect 2962 175879 3018 175888
rect 579526 168464 579582 168473
rect 579582 168422 579660 168450
rect 579526 168399 579582 168408
rect 579632 165889 579660 168422
rect 3054 165880 3110 165889
rect 3054 165815 3110 165824
rect 579618 165880 579674 165889
rect 579618 165815 579674 165824
rect 3068 162897 3096 165815
rect 3054 162888 3110 162897
rect 3054 162823 3110 162832
rect 579526 155544 579582 155553
rect 579582 155502 579660 155530
rect 579526 155479 579582 155488
rect 3054 153232 3110 153241
rect 3054 153167 3110 153176
rect 3068 149841 3096 153167
rect 579632 152697 579660 155502
rect 579618 152688 579674 152697
rect 579618 152623 579674 152632
rect 3054 149832 3110 149841
rect 3054 149767 3110 149776
rect 578790 142624 578846 142633
rect 578790 142559 578792 142568
rect 578844 142559 578846 142568
rect 580724 142588 580776 142594
rect 578792 142530 578844 142536
rect 580724 142530 580776 142536
rect 3054 140584 3110 140593
rect 3054 140519 3110 140528
rect 3068 136785 3096 140519
rect 580736 139369 580764 142530
rect 580722 139360 580778 139369
rect 580722 139295 580778 139304
rect 3054 136776 3110 136785
rect 3054 136711 3110 136720
rect 579526 129704 579582 129713
rect 579582 129662 579660 129690
rect 579526 129639 579582 129648
rect 3054 127936 3110 127945
rect 3054 127871 3110 127880
rect 3068 123729 3096 127871
rect 579632 126041 579660 129662
rect 579618 126032 579674 126041
rect 579618 125967 579674 125976
rect 3054 123720 3110 123729
rect 3054 123655 3110 123664
rect 578330 116784 578386 116793
rect 578330 116719 578332 116728
rect 578384 116719 578386 116728
rect 580264 116748 580316 116754
rect 578332 116690 578384 116696
rect 580264 116690 580316 116696
rect 2962 115288 3018 115297
rect 2962 115223 3018 115232
rect 2976 110673 3004 115223
rect 580276 112849 580304 116690
rect 580262 112840 580318 112849
rect 580262 112775 580318 112784
rect 2962 110664 3018 110673
rect 2962 110599 3018 110608
rect 579526 103864 579582 103873
rect 579526 103799 579582 103808
rect 579540 103514 579568 103799
rect 579540 103486 579844 103514
rect 3054 102640 3110 102649
rect 3054 102575 3110 102584
rect 3068 97617 3096 102575
rect 579816 99521 579844 103486
rect 579802 99512 579858 99521
rect 579802 99447 579858 99456
rect 3054 97608 3110 97617
rect 3054 97543 3110 97552
rect 579526 90944 579582 90953
rect 579582 90902 579660 90930
rect 579526 90879 579582 90888
rect 3054 89992 3110 90001
rect 3054 89927 3110 89936
rect 3068 84697 3096 89927
rect 579632 86193 579660 90902
rect 579618 86184 579674 86193
rect 579618 86119 579674 86128
rect 3054 84688 3110 84697
rect 3054 84623 3110 84632
rect 578882 78024 578938 78033
rect 578882 77959 578938 77968
rect 3422 77344 3478 77353
rect 3422 77279 3478 77288
rect 3436 71641 3464 77279
rect 578896 73001 578924 77959
rect 578882 72992 578938 73001
rect 578882 72927 578938 72936
rect 3422 71632 3478 71641
rect 3422 71567 3478 71576
rect 578238 65104 578294 65113
rect 578238 65039 578294 65048
rect 3054 64696 3110 64705
rect 3054 64631 3110 64640
rect 3068 58585 3096 64631
rect 578252 60722 578280 65039
rect 578240 60716 578292 60722
rect 578240 60658 578292 60664
rect 580816 60716 580868 60722
rect 580816 60658 580868 60664
rect 580828 59673 580856 60658
rect 580814 59664 580870 59673
rect 580814 59599 580870 59608
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 579526 52184 579582 52193
rect 579526 52119 579582 52128
rect 3422 52048 3478 52057
rect 3422 51983 3478 51992
rect 3436 45529 3464 51983
rect 579540 46345 579568 52119
rect 579526 46336 579582 46345
rect 579526 46271 579582 46280
rect 3422 45520 3478 45529
rect 3422 45455 3478 45464
rect 3422 39400 3478 39409
rect 3422 39335 3478 39344
rect 3436 32473 3464 39335
rect 578882 39264 578938 39273
rect 578882 39199 578938 39208
rect 578896 33153 578924 39199
rect 578882 33144 578938 33153
rect 578882 33079 578938 33088
rect 3422 32464 3478 32473
rect 3422 32399 3478 32408
rect 2962 26752 3018 26761
rect 2962 26687 3018 26696
rect 2976 19417 3004 26687
rect 578238 26344 578294 26353
rect 578238 26279 578294 26288
rect 578252 20670 578280 26279
rect 578240 20664 578292 20670
rect 578240 20606 578292 20612
rect 580632 20664 580684 20670
rect 580632 20606 580684 20612
rect 580644 19825 580672 20606
rect 580630 19816 580686 19825
rect 580630 19751 580686 19760
rect 2962 19408 3018 19417
rect 2962 19343 3018 19352
rect 3422 14104 3478 14113
rect 3422 14039 3478 14048
rect 3436 6497 3464 14039
rect 578882 13424 578938 13433
rect 578882 13359 578938 13368
rect 578896 6633 578924 13359
rect 578882 6624 578938 6633
rect 578882 6559 578938 6568
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 1676 4140 1728 4146
rect 1676 4082 1728 4088
rect 572 3800 624 3806
rect 572 3742 624 3748
rect 584 480 612 3742
rect 1688 480 1716 4082
rect 15936 4072 15988 4078
rect 15936 4014 15988 4020
rect 6460 4004 6512 4010
rect 6460 3946 6512 3952
rect 4068 3460 4120 3466
rect 4068 3402 4120 3408
rect 2872 3324 2924 3330
rect 2872 3266 2924 3272
rect 2884 480 2912 3266
rect 4080 480 4108 3402
rect 5262 3360 5318 3369
rect 5262 3295 5318 3304
rect 5276 480 5304 3295
rect 6472 480 6500 3946
rect 13544 3936 13596 3942
rect 13544 3878 13596 3884
rect 8760 3868 8812 3874
rect 8760 3810 8812 3816
rect 7656 3392 7708 3398
rect 7656 3334 7708 3340
rect 7668 480 7696 3334
rect 8772 480 8800 3810
rect 9956 3732 10008 3738
rect 9956 3674 10008 3680
rect 9968 480 9996 3674
rect 11152 3596 11204 3602
rect 11152 3538 11204 3544
rect 11164 480 11192 3538
rect 12348 3256 12400 3262
rect 12348 3198 12400 3204
rect 12360 480 12388 3198
rect 13556 480 13584 3878
rect 14740 3664 14792 3670
rect 14740 3606 14792 3612
rect 14752 480 14780 3606
rect 15948 480 15976 4014
rect 19168 3806 19196 6052
rect 20272 4146 20300 6052
rect 20260 4140 20312 4146
rect 20260 4082 20312 4088
rect 19156 3800 19208 3806
rect 19156 3742 19208 3748
rect 17040 3528 17092 3534
rect 17040 3470 17092 3476
rect 20626 3496 20682 3505
rect 17052 480 17080 3470
rect 20626 3431 20682 3440
rect 19432 3120 19484 3126
rect 19432 3062 19484 3068
rect 18236 3052 18288 3058
rect 18236 2994 18288 3000
rect 18248 480 18276 2994
rect 19444 480 19472 3062
rect 20640 480 20668 3431
rect 21376 3330 21404 6052
rect 21824 4140 21876 4146
rect 21824 4082 21876 4088
rect 21364 3324 21416 3330
rect 21364 3266 21416 3272
rect 21836 480 21864 4082
rect 22480 3466 22508 6052
rect 23020 3800 23072 3806
rect 23020 3742 23072 3748
rect 22468 3460 22520 3466
rect 22468 3402 22520 3408
rect 23032 480 23060 3742
rect 23584 3369 23612 6052
rect 24688 4010 24716 6052
rect 24676 4004 24728 4010
rect 24676 3946 24728 3952
rect 25792 3398 25820 6052
rect 26896 3874 26924 6052
rect 26884 3868 26936 3874
rect 26884 3810 26936 3816
rect 28000 3738 28028 6052
rect 27988 3732 28040 3738
rect 27988 3674 28040 3680
rect 29104 3602 29132 6052
rect 29092 3596 29144 3602
rect 29092 3538 29144 3544
rect 30104 3460 30156 3466
rect 30104 3402 30156 3408
rect 25780 3392 25832 3398
rect 23570 3360 23626 3369
rect 25780 3334 25832 3340
rect 28906 3360 28962 3369
rect 23570 3295 23626 3304
rect 26516 3324 26568 3330
rect 28906 3295 28962 3304
rect 26516 3266 26568 3272
rect 24216 3188 24268 3194
rect 24216 3130 24268 3136
rect 24228 480 24256 3130
rect 25320 2984 25372 2990
rect 25320 2926 25372 2932
rect 25332 480 25360 2926
rect 26528 480 26556 3266
rect 27712 2916 27764 2922
rect 27712 2858 27764 2864
rect 27724 480 27752 2858
rect 28920 480 28948 3295
rect 30116 480 30144 3402
rect 30208 3262 30236 6052
rect 31312 3942 31340 6052
rect 31300 3936 31352 3942
rect 31300 3878 31352 3884
rect 31300 3732 31352 3738
rect 31300 3674 31352 3680
rect 30196 3256 30248 3262
rect 30196 3198 30248 3204
rect 31312 480 31340 3674
rect 32416 3670 32444 6052
rect 33520 4078 33548 6052
rect 33508 4072 33560 4078
rect 33508 4014 33560 4020
rect 32496 3868 32548 3874
rect 32496 3810 32548 3816
rect 32404 3664 32456 3670
rect 32404 3606 32456 3612
rect 32508 1986 32536 3810
rect 34624 3534 34652 6052
rect 34796 3664 34848 3670
rect 34796 3606 34848 3612
rect 34612 3528 34664 3534
rect 34612 3470 34664 3476
rect 33600 3392 33652 3398
rect 33600 3334 33652 3340
rect 32416 1958 32536 1986
rect 32416 480 32444 1958
rect 33612 480 33640 3334
rect 34808 480 34836 3606
rect 35728 3058 35756 6052
rect 36832 3126 36860 6052
rect 37936 3505 37964 6052
rect 39040 4146 39068 6052
rect 39028 4140 39080 4146
rect 39028 4082 39080 4088
rect 39580 4004 39632 4010
rect 39580 3946 39632 3952
rect 38384 3936 38436 3942
rect 38384 3878 38436 3884
rect 37922 3496 37978 3505
rect 37922 3431 37978 3440
rect 37188 3256 37240 3262
rect 37188 3198 37240 3204
rect 36820 3120 36872 3126
rect 36820 3062 36872 3068
rect 35716 3052 35768 3058
rect 35716 2994 35768 3000
rect 35992 2848 36044 2854
rect 35992 2790 36044 2796
rect 36004 480 36032 2790
rect 37200 480 37228 3198
rect 38396 480 38424 3878
rect 39592 480 39620 3946
rect 40144 3806 40172 6052
rect 40684 4072 40736 4078
rect 40684 4014 40736 4020
rect 40132 3800 40184 3806
rect 40132 3742 40184 3748
rect 40696 480 40724 4014
rect 41248 3194 41276 6052
rect 41880 3800 41932 3806
rect 41880 3742 41932 3748
rect 41236 3188 41288 3194
rect 41236 3130 41288 3136
rect 41892 480 41920 3742
rect 42352 2990 42380 6052
rect 43076 4140 43128 4146
rect 43076 4082 43128 4088
rect 42340 2984 42392 2990
rect 42340 2926 42392 2932
rect 43088 480 43116 4082
rect 43456 3330 43484 6052
rect 43444 3324 43496 3330
rect 43444 3266 43496 3272
rect 44272 3120 44324 3126
rect 44272 3062 44324 3068
rect 44284 480 44312 3062
rect 44560 2922 44588 6052
rect 45468 3528 45520 3534
rect 45468 3470 45520 3476
rect 44548 2916 44600 2922
rect 44548 2858 44600 2864
rect 45480 480 45508 3470
rect 45664 3369 45692 6052
rect 46664 3596 46716 3602
rect 46664 3538 46716 3544
rect 45650 3360 45706 3369
rect 45650 3295 45706 3304
rect 46676 480 46704 3538
rect 46768 3466 46796 6052
rect 47872 3738 47900 6052
rect 48976 3874 49004 6052
rect 48964 3868 49016 3874
rect 48964 3810 49016 3816
rect 47860 3732 47912 3738
rect 47860 3674 47912 3680
rect 46756 3460 46808 3466
rect 46756 3402 46808 3408
rect 48964 3460 49016 3466
rect 48964 3402 49016 3408
rect 47860 3188 47912 3194
rect 47860 3130 47912 3136
rect 47872 480 47900 3130
rect 48976 480 49004 3402
rect 50080 3398 50108 6052
rect 50160 3732 50212 3738
rect 50160 3674 50212 3680
rect 50068 3392 50120 3398
rect 50068 3334 50120 3340
rect 50172 480 50200 3674
rect 51184 3670 51212 6052
rect 51172 3664 51224 3670
rect 51172 3606 51224 3612
rect 51356 3392 51408 3398
rect 51356 3334 51408 3340
rect 51368 480 51396 3334
rect 52288 2854 52316 6052
rect 53392 3330 53420 6052
rect 54496 3942 54524 6052
rect 55600 4010 55628 6052
rect 56704 4078 56732 6052
rect 56692 4072 56744 4078
rect 56692 4014 56744 4020
rect 55588 4004 55640 4010
rect 55588 3946 55640 3952
rect 54484 3936 54536 3942
rect 54484 3878 54536 3884
rect 57244 3936 57296 3942
rect 57244 3878 57296 3884
rect 53748 3868 53800 3874
rect 53748 3810 53800 3816
rect 53380 3324 53432 3330
rect 53380 3266 53432 3272
rect 52552 3256 52604 3262
rect 52552 3198 52604 3204
rect 52276 2848 52328 2854
rect 52276 2790 52328 2796
rect 52564 480 52592 3198
rect 53760 480 53788 3810
rect 56048 3664 56100 3670
rect 56048 3606 56100 3612
rect 54944 3324 54996 3330
rect 54944 3266 54996 3272
rect 54956 480 54984 3266
rect 56060 480 56088 3606
rect 57256 480 57284 3878
rect 57808 3806 57836 6052
rect 58912 4146 58940 6052
rect 58900 4140 58952 4146
rect 58900 4082 58952 4088
rect 58440 4004 58492 4010
rect 58440 3946 58492 3952
rect 57796 3800 57848 3806
rect 57796 3742 57848 3748
rect 58452 480 58480 3946
rect 60016 3126 60044 6052
rect 61120 3534 61148 6052
rect 62028 4072 62080 4078
rect 62028 4014 62080 4020
rect 61108 3528 61160 3534
rect 61108 3470 61160 3476
rect 60004 3120 60056 3126
rect 60004 3062 60056 3068
rect 60832 3120 60884 3126
rect 60832 3062 60884 3068
rect 59636 2984 59688 2990
rect 59636 2926 59688 2932
rect 59648 480 59676 2926
rect 60844 480 60872 3062
rect 62040 480 62068 4014
rect 62224 3602 62252 6052
rect 63224 3800 63276 3806
rect 63224 3742 63276 3748
rect 62212 3596 62264 3602
rect 62212 3538 62264 3544
rect 63236 480 63264 3742
rect 63328 3194 63356 6052
rect 64328 3596 64380 3602
rect 64328 3538 64380 3544
rect 63316 3188 63368 3194
rect 63316 3130 63368 3136
rect 64340 480 64368 3538
rect 64432 3466 64460 6052
rect 65536 3738 65564 6052
rect 65524 3732 65576 3738
rect 65524 3674 65576 3680
rect 64420 3460 64472 3466
rect 64420 3402 64472 3408
rect 66640 3398 66668 6052
rect 66720 4140 66772 4146
rect 66720 4082 66772 4088
rect 66628 3392 66680 3398
rect 66628 3334 66680 3340
rect 65524 3188 65576 3194
rect 65524 3130 65576 3136
rect 65536 480 65564 3130
rect 66732 480 66760 4082
rect 67744 3262 67772 6052
rect 68848 3874 68876 6052
rect 68836 3868 68888 3874
rect 68836 3810 68888 3816
rect 67916 3528 67968 3534
rect 67916 3470 67968 3476
rect 67732 3256 67784 3262
rect 67732 3198 67784 3204
rect 67928 480 67956 3470
rect 69952 3330 69980 6052
rect 71056 3670 71084 6052
rect 72160 3942 72188 6052
rect 73264 4010 73292 6052
rect 73252 4004 73304 4010
rect 73252 3946 73304 3952
rect 72148 3936 72200 3942
rect 72148 3878 72200 3884
rect 71504 3868 71556 3874
rect 71504 3810 71556 3816
rect 71044 3664 71096 3670
rect 71044 3606 71096 3612
rect 70308 3460 70360 3466
rect 70308 3402 70360 3408
rect 69940 3324 69992 3330
rect 69940 3266 69992 3272
rect 69112 3052 69164 3058
rect 69112 2994 69164 3000
rect 69124 480 69152 2994
rect 70320 480 70348 3402
rect 71516 480 71544 3810
rect 73804 3324 73856 3330
rect 73804 3266 73856 3272
rect 72608 3256 72660 3262
rect 72608 3198 72660 3204
rect 72620 480 72648 3198
rect 73816 480 73844 3266
rect 74368 2990 74396 6052
rect 75000 3732 75052 3738
rect 75000 3674 75052 3680
rect 74356 2984 74408 2990
rect 74356 2926 74408 2932
rect 75012 480 75040 3674
rect 75472 3126 75500 6052
rect 76576 4078 76604 6052
rect 76564 4072 76616 4078
rect 76564 4014 76616 4020
rect 77392 4072 77444 4078
rect 77392 4014 77444 4020
rect 76196 3392 76248 3398
rect 76196 3334 76248 3340
rect 75460 3120 75512 3126
rect 75460 3062 75512 3068
rect 76208 480 76236 3334
rect 77404 480 77432 4014
rect 77680 3806 77708 6052
rect 78588 3936 78640 3942
rect 78588 3878 78640 3884
rect 77668 3800 77720 3806
rect 77668 3742 77720 3748
rect 78600 480 78628 3878
rect 78784 3602 78812 6052
rect 79692 3800 79744 3806
rect 79692 3742 79744 3748
rect 78772 3596 78824 3602
rect 78772 3538 78824 3544
rect 79704 480 79732 3742
rect 79888 3194 79916 6052
rect 80992 4146 81020 6052
rect 81728 6038 82110 6066
rect 80980 4140 81032 4146
rect 80980 4082 81032 4088
rect 80888 3596 80940 3602
rect 80888 3538 80940 3544
rect 79876 3188 79928 3194
rect 79876 3130 79928 3136
rect 80900 480 80928 3538
rect 81728 3534 81756 6038
rect 82084 3664 82136 3670
rect 82084 3606 82136 3612
rect 81716 3528 81768 3534
rect 81716 3470 81768 3476
rect 82096 480 82124 3606
rect 83200 3058 83228 6052
rect 83280 4140 83332 4146
rect 83280 4082 83332 4088
rect 83188 3052 83240 3058
rect 83188 2994 83240 3000
rect 83292 480 83320 4082
rect 84304 3466 84332 6052
rect 84476 4004 84528 4010
rect 84476 3946 84528 3952
rect 84292 3460 84344 3466
rect 84292 3402 84344 3408
rect 84488 480 84516 3946
rect 85408 3874 85436 6052
rect 85396 3868 85448 3874
rect 85396 3810 85448 3816
rect 86512 3262 86540 6052
rect 86868 3528 86920 3534
rect 86868 3470 86920 3476
rect 86500 3256 86552 3262
rect 86500 3198 86552 3204
rect 85672 3188 85724 3194
rect 85672 3130 85724 3136
rect 85684 480 85712 3130
rect 86880 480 86908 3470
rect 87616 3330 87644 6052
rect 88720 3738 88748 6052
rect 89168 3868 89220 3874
rect 89168 3810 89220 3816
rect 88708 3732 88760 3738
rect 88708 3674 88760 3680
rect 87972 3460 88024 3466
rect 87972 3402 88024 3408
rect 87604 3324 87656 3330
rect 87604 3266 87656 3272
rect 87984 480 88012 3402
rect 89180 480 89208 3810
rect 89824 3398 89852 6052
rect 90928 4078 90956 6052
rect 90916 4072 90968 4078
rect 90916 4014 90968 4020
rect 92032 3942 92060 6052
rect 92020 3936 92072 3942
rect 92020 3878 92072 3884
rect 92756 3936 92808 3942
rect 92756 3878 92808 3884
rect 91560 3732 91612 3738
rect 91560 3674 91612 3680
rect 89812 3392 89864 3398
rect 89812 3334 89864 3340
rect 90364 3256 90416 3262
rect 90364 3198 90416 3204
rect 90376 480 90404 3198
rect 91572 480 91600 3674
rect 92768 480 92796 3878
rect 93136 3806 93164 6052
rect 93952 4072 94004 4078
rect 93952 4014 94004 4020
rect 93124 3800 93176 3806
rect 93124 3742 93176 3748
rect 93964 480 93992 4014
rect 94240 3602 94268 6052
rect 95344 3670 95372 6052
rect 96448 4146 96476 6052
rect 96436 4140 96488 4146
rect 96436 4082 96488 4088
rect 97448 4140 97500 4146
rect 97448 4082 97500 4088
rect 96252 3800 96304 3806
rect 96252 3742 96304 3748
rect 95332 3664 95384 3670
rect 95332 3606 95384 3612
rect 94228 3596 94280 3602
rect 94228 3538 94280 3544
rect 95148 3392 95200 3398
rect 95148 3334 95200 3340
rect 95160 480 95188 3334
rect 96264 480 96292 3742
rect 97460 480 97488 4082
rect 97552 4010 97580 6052
rect 98288 6038 98670 6066
rect 97540 4004 97592 4010
rect 97540 3946 97592 3952
rect 98288 3194 98316 6038
rect 98644 3596 98696 3602
rect 98644 3538 98696 3544
rect 98276 3188 98328 3194
rect 98276 3130 98328 3136
rect 98656 480 98684 3538
rect 99760 3534 99788 6052
rect 99840 3664 99892 3670
rect 99840 3606 99892 3612
rect 99748 3528 99800 3534
rect 99748 3470 99800 3476
rect 99852 480 99880 3606
rect 100864 3466 100892 6052
rect 101036 4004 101088 4010
rect 101036 3946 101088 3952
rect 100852 3460 100904 3466
rect 100852 3402 100904 3408
rect 101048 480 101076 3946
rect 101968 3874 101996 6052
rect 101956 3868 102008 3874
rect 101956 3810 102008 3816
rect 103072 3262 103100 6052
rect 103336 3868 103388 3874
rect 103336 3810 103388 3816
rect 103060 3256 103112 3262
rect 103060 3198 103112 3204
rect 102232 3120 102284 3126
rect 102232 3062 102284 3068
rect 102244 480 102272 3062
rect 103348 480 103376 3810
rect 104176 3738 104204 6052
rect 105280 3942 105308 6052
rect 106384 4078 106412 6052
rect 106372 4072 106424 4078
rect 106372 4014 106424 4020
rect 105268 3936 105320 3942
rect 105268 3878 105320 3884
rect 104164 3732 104216 3738
rect 104164 3674 104216 3680
rect 105728 3528 105780 3534
rect 105728 3470 105780 3476
rect 104532 3460 104584 3466
rect 104532 3402 104584 3408
rect 104544 480 104572 3402
rect 105740 480 105768 3470
rect 107488 3398 107516 6052
rect 108120 3936 108172 3942
rect 108120 3878 108172 3884
rect 107476 3392 107528 3398
rect 107476 3334 107528 3340
rect 106924 3256 106976 3262
rect 106924 3198 106976 3204
rect 106936 480 106964 3198
rect 108132 480 108160 3878
rect 108592 3806 108620 6052
rect 109696 4146 109724 6052
rect 109684 4140 109736 4146
rect 109684 4082 109736 4088
rect 108580 3800 108632 3806
rect 108580 3742 108632 3748
rect 110512 3800 110564 3806
rect 110512 3742 110564 3748
rect 109316 3324 109368 3330
rect 109316 3266 109368 3272
rect 109328 480 109356 3266
rect 110524 480 110552 3742
rect 110800 3602 110828 6052
rect 111904 3670 111932 6052
rect 112812 4140 112864 4146
rect 112812 4082 112864 4088
rect 111892 3664 111944 3670
rect 111892 3606 111944 3612
rect 110788 3596 110840 3602
rect 110788 3538 110840 3544
rect 111616 3596 111668 3602
rect 111616 3538 111668 3544
rect 111628 480 111656 3538
rect 112824 480 112852 4082
rect 113008 4010 113036 6052
rect 112996 4004 113048 4010
rect 112996 3946 113048 3952
rect 114008 3664 114060 3670
rect 114008 3606 114060 3612
rect 114020 480 114048 3606
rect 114112 3126 114140 6052
rect 115216 3874 115244 6052
rect 115296 4004 115348 4010
rect 115296 3946 115348 3952
rect 115204 3868 115256 3874
rect 115204 3810 115256 3816
rect 114100 3120 114152 3126
rect 114100 3062 114152 3068
rect 115308 1986 115336 3946
rect 116320 3466 116348 6052
rect 116400 3868 116452 3874
rect 116400 3810 116452 3816
rect 116308 3460 116360 3466
rect 116308 3402 116360 3408
rect 115216 1958 115336 1986
rect 115216 480 115244 1958
rect 116412 480 116440 3810
rect 117424 3534 117452 6052
rect 117596 3732 117648 3738
rect 117596 3674 117648 3680
rect 117412 3528 117464 3534
rect 117412 3470 117464 3476
rect 117608 480 117636 3674
rect 118528 3262 118556 6052
rect 119632 3942 119660 6052
rect 119896 4072 119948 4078
rect 119896 4014 119948 4020
rect 119620 3936 119672 3942
rect 119620 3878 119672 3884
rect 118792 3392 118844 3398
rect 118792 3334 118844 3340
rect 118516 3256 118568 3262
rect 118516 3198 118568 3204
rect 118804 480 118832 3334
rect 119908 480 119936 4014
rect 120736 3330 120764 6052
rect 121840 3806 121868 6052
rect 122288 3936 122340 3942
rect 122288 3878 122340 3884
rect 121828 3800 121880 3806
rect 121828 3742 121880 3748
rect 121092 3460 121144 3466
rect 121092 3402 121144 3408
rect 120724 3324 120776 3330
rect 120724 3266 120776 3272
rect 121104 480 121132 3402
rect 122300 480 122328 3878
rect 122944 3602 122972 6052
rect 124048 4146 124076 6052
rect 124036 4140 124088 4146
rect 124036 4082 124088 4088
rect 124680 4140 124732 4146
rect 124680 4082 124732 4088
rect 123484 3800 123536 3806
rect 123484 3742 123536 3748
rect 122932 3596 122984 3602
rect 122932 3538 122984 3544
rect 123496 480 123524 3742
rect 124692 480 124720 4082
rect 125152 3670 125180 6052
rect 126256 4010 126284 6052
rect 126244 4004 126296 4010
rect 126244 3946 126296 3952
rect 126980 4004 127032 4010
rect 126980 3946 127032 3952
rect 125140 3664 125192 3670
rect 125140 3606 125192 3612
rect 125876 3324 125928 3330
rect 125876 3266 125928 3272
rect 125888 480 125916 3266
rect 126992 480 127020 3946
rect 127360 3874 127388 6052
rect 127348 3868 127400 3874
rect 127348 3810 127400 3816
rect 128464 3738 128492 6052
rect 128452 3732 128504 3738
rect 128452 3674 128504 3680
rect 128176 3596 128228 3602
rect 128176 3538 128228 3544
rect 128188 480 128216 3538
rect 129372 3528 129424 3534
rect 129372 3470 129424 3476
rect 129384 480 129412 3470
rect 129568 3398 129596 6052
rect 130672 4078 130700 6052
rect 131408 6038 131790 6066
rect 130660 4072 130712 4078
rect 130660 4014 130712 4020
rect 131408 3466 131436 6038
rect 132880 3942 132908 6052
rect 132960 4072 133012 4078
rect 132960 4014 133012 4020
rect 132868 3936 132920 3942
rect 132868 3878 132920 3884
rect 131764 3664 131816 3670
rect 131764 3606 131816 3612
rect 131396 3460 131448 3466
rect 131396 3402 131448 3408
rect 129556 3392 129608 3398
rect 129556 3334 129608 3340
rect 130568 3392 130620 3398
rect 130568 3334 130620 3340
rect 130580 480 130608 3334
rect 131776 480 131804 3606
rect 132972 480 133000 4014
rect 133984 3806 134012 6052
rect 135088 4146 135116 6052
rect 135076 4140 135128 4146
rect 135076 4082 135128 4088
rect 134156 3936 134208 3942
rect 134156 3878 134208 3884
rect 133972 3800 134024 3806
rect 133972 3742 134024 3748
rect 134168 480 134196 3878
rect 135260 3460 135312 3466
rect 135260 3402 135312 3408
rect 135272 480 135300 3402
rect 136192 3330 136220 6052
rect 136456 4140 136508 4146
rect 136456 4082 136508 4088
rect 136180 3324 136232 3330
rect 136180 3266 136232 3272
rect 136468 480 136496 4082
rect 137296 4010 137324 6052
rect 137284 4004 137336 4010
rect 137284 3946 137336 3952
rect 137652 3868 137704 3874
rect 137652 3810 137704 3816
rect 137664 480 137692 3810
rect 138400 3602 138428 6052
rect 138848 3732 138900 3738
rect 138848 3674 138900 3680
rect 138388 3596 138440 3602
rect 138388 3538 138440 3544
rect 138860 480 138888 3674
rect 139504 3534 139532 6052
rect 140044 3800 140096 3806
rect 140044 3742 140096 3748
rect 139492 3528 139544 3534
rect 139492 3470 139544 3476
rect 140056 480 140084 3742
rect 140608 3398 140636 6052
rect 141712 3670 141740 6052
rect 142816 4078 142844 6052
rect 142804 4072 142856 4078
rect 142804 4014 142856 4020
rect 143540 4072 143592 4078
rect 143540 4014 143592 4020
rect 141700 3664 141752 3670
rect 141700 3606 141752 3612
rect 141240 3528 141292 3534
rect 141240 3470 141292 3476
rect 140596 3392 140648 3398
rect 140596 3334 140648 3340
rect 141252 480 141280 3470
rect 142436 3052 142488 3058
rect 142436 2994 142488 3000
rect 142448 480 142476 2994
rect 143552 480 143580 4014
rect 143920 3942 143948 6052
rect 143908 3936 143960 3942
rect 143908 3878 143960 3884
rect 144736 3664 144788 3670
rect 144736 3606 144788 3612
rect 144748 480 144776 3606
rect 145024 3466 145052 6052
rect 146128 4146 146156 6052
rect 146116 4140 146168 4146
rect 146116 4082 146168 4088
rect 147232 3874 147260 6052
rect 147968 6038 148350 6066
rect 147220 3868 147272 3874
rect 147220 3810 147272 3816
rect 147968 3738 147996 6038
rect 148324 3868 148376 3874
rect 148324 3810 148376 3816
rect 147956 3732 148008 3738
rect 147956 3674 148008 3680
rect 145932 3596 145984 3602
rect 145932 3538 145984 3544
rect 145012 3460 145064 3466
rect 145012 3402 145064 3408
rect 145944 480 145972 3538
rect 147128 3460 147180 3466
rect 147128 3402 147180 3408
rect 147140 480 147168 3402
rect 148336 480 148364 3810
rect 149440 3806 149468 6052
rect 149520 3936 149572 3942
rect 149520 3878 149572 3884
rect 149428 3800 149480 3806
rect 149428 3742 149480 3748
rect 149532 480 149560 3878
rect 150544 3534 150572 6052
rect 150624 4004 150676 4010
rect 150624 3946 150676 3952
rect 150532 3528 150584 3534
rect 150532 3470 150584 3476
rect 150636 480 150664 3946
rect 151648 3058 151676 6052
rect 152752 4078 152780 6052
rect 152740 4072 152792 4078
rect 152740 4014 152792 4020
rect 153856 3670 153884 6052
rect 154212 4072 154264 4078
rect 154212 4014 154264 4020
rect 153844 3664 153896 3670
rect 153844 3606 153896 3612
rect 153016 3528 153068 3534
rect 153016 3470 153068 3476
rect 151636 3052 151688 3058
rect 151636 2994 151688 3000
rect 151820 3052 151872 3058
rect 151820 2994 151872 3000
rect 151832 480 151860 2994
rect 153028 480 153056 3470
rect 154224 480 154252 4014
rect 154960 3602 154988 6052
rect 154948 3596 155000 3602
rect 154948 3538 155000 3544
rect 156064 3466 156092 6052
rect 157168 3874 157196 6052
rect 157800 4140 157852 4146
rect 157800 4082 157852 4088
rect 157156 3868 157208 3874
rect 157156 3810 157208 3816
rect 156604 3596 156656 3602
rect 156604 3538 156656 3544
rect 156052 3460 156104 3466
rect 156052 3402 156104 3408
rect 155408 2916 155460 2922
rect 155408 2858 155460 2864
rect 155420 480 155448 2858
rect 156616 480 156644 3538
rect 157812 480 157840 4082
rect 158272 3942 158300 6052
rect 159376 4010 159404 6052
rect 159364 4004 159416 4010
rect 159364 3946 159416 3952
rect 158260 3936 158312 3942
rect 158260 3878 158312 3884
rect 160100 3936 160152 3942
rect 160100 3878 160152 3884
rect 158904 3460 158956 3466
rect 158904 3402 158956 3408
rect 158916 480 158944 3402
rect 160112 480 160140 3878
rect 160480 3058 160508 6052
rect 161296 3868 161348 3874
rect 161296 3810 161348 3816
rect 160468 3052 160520 3058
rect 160468 2994 160520 3000
rect 161308 480 161336 3810
rect 161584 3534 161612 6052
rect 162688 4078 162716 6052
rect 162676 4072 162728 4078
rect 162676 4014 162728 4020
rect 161572 3528 161624 3534
rect 161572 3470 161624 3476
rect 163688 3528 163740 3534
rect 163688 3470 163740 3476
rect 162492 2984 162544 2990
rect 162492 2926 162544 2932
rect 162504 480 162532 2926
rect 163700 480 163728 3470
rect 163792 2922 163820 6052
rect 164896 3602 164924 6052
rect 166000 4146 166028 6052
rect 165988 4140 166040 4146
rect 165988 4082 166040 4088
rect 164884 3596 164936 3602
rect 164884 3538 164936 3544
rect 167104 3466 167132 6052
rect 168208 3942 168236 6052
rect 168380 4072 168432 4078
rect 168380 4014 168432 4020
rect 168196 3936 168248 3942
rect 168196 3878 168248 3884
rect 167184 3800 167236 3806
rect 167184 3742 167236 3748
rect 167092 3460 167144 3466
rect 167092 3402 167144 3408
rect 164884 3120 164936 3126
rect 164884 3062 164936 3068
rect 163780 2916 163832 2922
rect 163780 2858 163832 2864
rect 164896 480 164924 3062
rect 166080 3052 166132 3058
rect 166080 2994 166132 3000
rect 166092 480 166120 2994
rect 167196 480 167224 3742
rect 168392 480 168420 4014
rect 169312 3874 169340 6052
rect 169300 3868 169352 3874
rect 169300 3810 169352 3816
rect 169576 3596 169628 3602
rect 169576 3538 169628 3544
rect 169588 480 169616 3538
rect 170416 2990 170444 6052
rect 171520 3534 171548 6052
rect 171508 3528 171560 3534
rect 171508 3470 171560 3476
rect 170772 3460 170824 3466
rect 170772 3402 170824 3408
rect 170404 2984 170456 2990
rect 170404 2926 170456 2932
rect 170784 480 170812 3402
rect 172624 3126 172652 6052
rect 172612 3120 172664 3126
rect 172612 3062 172664 3068
rect 173728 3058 173756 6052
rect 174268 4140 174320 4146
rect 174268 4082 174320 4088
rect 173716 3052 173768 3058
rect 173716 2994 173768 3000
rect 171968 2984 172020 2990
rect 171968 2926 172020 2932
rect 171980 480 172008 2926
rect 173164 2916 173216 2922
rect 173164 2858 173216 2864
rect 173176 480 173204 2858
rect 174280 480 174308 4082
rect 174832 3806 174860 6052
rect 175936 4078 175964 6052
rect 175924 4072 175976 4078
rect 175924 4014 175976 4020
rect 176660 4072 176712 4078
rect 176660 4014 176712 4020
rect 174820 3800 174872 3806
rect 174820 3742 174872 3748
rect 175464 3800 175516 3806
rect 175464 3742 175516 3748
rect 175476 480 175504 3742
rect 176672 480 176700 4014
rect 177040 3602 177068 6052
rect 177856 3732 177908 3738
rect 177856 3674 177908 3680
rect 177028 3596 177080 3602
rect 177028 3538 177080 3544
rect 177868 480 177896 3674
rect 178144 3466 178172 6052
rect 179052 3936 179104 3942
rect 179052 3878 179104 3884
rect 178132 3460 178184 3466
rect 178132 3402 178184 3408
rect 179064 480 179092 3878
rect 179248 2990 179276 6052
rect 180248 4004 180300 4010
rect 180248 3946 180300 3952
rect 179236 2984 179288 2990
rect 179236 2926 179288 2932
rect 180260 480 180288 3946
rect 180352 2922 180380 6052
rect 181456 4146 181484 6052
rect 181444 4140 181496 4146
rect 181444 4082 181496 4088
rect 182560 3806 182588 6052
rect 183664 4078 183692 6052
rect 183652 4072 183704 4078
rect 183652 4014 183704 4020
rect 182548 3800 182600 3806
rect 182548 3742 182600 3748
rect 184768 3738 184796 6052
rect 185872 3942 185900 6052
rect 186976 4010 187004 6052
rect 186964 4004 187016 4010
rect 186964 3946 187016 3952
rect 185860 3936 185912 3942
rect 185860 3878 185912 3884
rect 184756 3732 184808 3738
rect 184756 3674 184808 3680
rect 187332 3528 187384 3534
rect 187332 3470 187384 3476
rect 181444 3256 181496 3262
rect 181444 3198 181496 3204
rect 180340 2916 180392 2922
rect 180340 2858 180392 2864
rect 181456 480 181484 3198
rect 182548 3188 182600 3194
rect 182548 3130 182600 3136
rect 182560 480 182588 3130
rect 184940 3120 184992 3126
rect 184940 3062 184992 3068
rect 183744 2984 183796 2990
rect 183744 2926 183796 2932
rect 183756 480 183784 2926
rect 184952 480 184980 3062
rect 186136 3052 186188 3058
rect 186136 2994 186188 3000
rect 186148 480 186176 2994
rect 187344 480 187372 3470
rect 188080 3262 188108 6052
rect 188528 3460 188580 3466
rect 188528 3402 188580 3408
rect 188068 3256 188120 3262
rect 188068 3198 188120 3204
rect 188540 480 188568 3402
rect 189184 3194 189212 6052
rect 189724 4004 189776 4010
rect 189724 3946 189776 3952
rect 189172 3188 189224 3194
rect 189172 3130 189224 3136
rect 189736 480 189764 3946
rect 190288 2990 190316 6052
rect 191392 3126 191420 6052
rect 192024 3188 192076 3194
rect 192024 3130 192076 3136
rect 191380 3120 191432 3126
rect 191380 3062 191432 3068
rect 190276 2984 190328 2990
rect 190276 2926 190328 2932
rect 190828 2916 190880 2922
rect 190828 2858 190880 2864
rect 190840 480 190868 2858
rect 192036 480 192064 3130
rect 192496 3058 192524 6052
rect 193220 3596 193272 3602
rect 193220 3538 193272 3544
rect 192484 3052 192536 3058
rect 192484 2994 192536 3000
rect 193232 480 193260 3538
rect 193600 3534 193628 6052
rect 193588 3528 193640 3534
rect 193588 3470 193640 3476
rect 194704 3466 194732 6052
rect 195808 4010 195836 6052
rect 195796 4004 195848 4010
rect 195796 3946 195848 3952
rect 194692 3460 194744 3466
rect 194692 3402 194744 3408
rect 195612 3120 195664 3126
rect 195612 3062 195664 3068
rect 194416 2984 194468 2990
rect 194416 2926 194468 2932
rect 194428 480 194456 2926
rect 195624 480 195652 3062
rect 196808 3052 196860 3058
rect 196808 2994 196860 3000
rect 196820 480 196848 2994
rect 196912 2922 196940 6052
rect 197912 3800 197964 3806
rect 197912 3742 197964 3748
rect 196900 2916 196952 2922
rect 196900 2858 196952 2864
rect 197924 480 197952 3742
rect 198016 3194 198044 6052
rect 199120 3602 199148 6052
rect 199108 3596 199160 3602
rect 199108 3538 199160 3544
rect 199108 3460 199160 3466
rect 199108 3402 199160 3408
rect 198004 3188 198056 3194
rect 198004 3130 198056 3136
rect 199120 480 199148 3402
rect 200224 2990 200252 6052
rect 201328 3126 201356 6052
rect 201500 3256 201552 3262
rect 201500 3198 201552 3204
rect 201316 3120 201368 3126
rect 201316 3062 201368 3068
rect 200212 2984 200264 2990
rect 200212 2926 200264 2932
rect 200304 2984 200356 2990
rect 200304 2926 200356 2932
rect 200316 480 200344 2926
rect 201512 480 201540 3198
rect 202432 3058 202460 6052
rect 203536 3806 203564 6052
rect 203524 3800 203576 3806
rect 203524 3742 203576 3748
rect 204640 3466 204668 6052
rect 204628 3460 204680 3466
rect 204628 3402 204680 3408
rect 203892 3188 203944 3194
rect 203892 3130 203944 3136
rect 202420 3052 202472 3058
rect 202420 2994 202472 3000
rect 202696 2916 202748 2922
rect 202696 2858 202748 2864
rect 202708 480 202736 2858
rect 203904 480 203932 3130
rect 205088 3120 205140 3126
rect 205088 3062 205140 3068
rect 205100 480 205128 3062
rect 205744 2990 205772 6052
rect 206848 3262 206876 6052
rect 206836 3256 206888 3262
rect 206836 3198 206888 3204
rect 207388 3052 207440 3058
rect 207388 2994 207440 3000
rect 205732 2984 205784 2990
rect 205732 2926 205784 2932
rect 206192 2984 206244 2990
rect 206192 2926 206244 2932
rect 206204 480 206232 2926
rect 207400 480 207428 2994
rect 207952 2922 207980 6052
rect 208584 3800 208636 3806
rect 208584 3742 208636 3748
rect 207940 2916 207992 2922
rect 207940 2858 207992 2864
rect 208596 480 208624 3742
rect 209056 3194 209084 6052
rect 209044 3188 209096 3194
rect 209044 3130 209096 3136
rect 210160 3126 210188 6052
rect 210976 3256 211028 3262
rect 210976 3198 211028 3204
rect 210148 3120 210200 3126
rect 210148 3062 210200 3068
rect 209780 2848 209832 2854
rect 209780 2790 209832 2796
rect 209792 480 209820 2790
rect 210988 480 211016 3198
rect 211264 2990 211292 6052
rect 212368 3058 212396 6052
rect 213472 3806 213500 6052
rect 213460 3800 213512 3806
rect 213460 3742 213512 3748
rect 213368 3188 213420 3194
rect 213368 3130 213420 3136
rect 212356 3052 212408 3058
rect 212356 2994 212408 3000
rect 211252 2984 211304 2990
rect 211252 2926 211304 2932
rect 212172 2916 212224 2922
rect 212172 2858 212224 2864
rect 212184 480 212212 2858
rect 213380 480 213408 3130
rect 214472 2984 214524 2990
rect 214472 2926 214524 2932
rect 214484 480 214512 2926
rect 214576 2854 214604 6052
rect 215680 3262 215708 6052
rect 215668 3256 215720 3262
rect 215668 3198 215720 3204
rect 215668 3120 215720 3126
rect 215668 3062 215720 3068
rect 214564 2848 214616 2854
rect 214564 2790 214616 2796
rect 215680 480 215708 3062
rect 216784 2922 216812 6052
rect 217888 3194 217916 6052
rect 218060 3800 218112 3806
rect 218060 3742 218112 3748
rect 217876 3188 217928 3194
rect 217876 3130 217928 3136
rect 216864 3052 216916 3058
rect 216864 2994 216916 3000
rect 216772 2916 216824 2922
rect 216772 2858 216824 2864
rect 216876 480 216904 2994
rect 218072 480 218100 3742
rect 218992 2990 219020 6052
rect 219256 3528 219308 3534
rect 219256 3470 219308 3476
rect 218980 2984 219032 2990
rect 218980 2926 219032 2932
rect 219268 480 219296 3470
rect 220096 3126 220124 6052
rect 220084 3120 220136 3126
rect 220084 3062 220136 3068
rect 221200 3058 221228 6052
rect 222304 3806 222332 6052
rect 222292 3800 222344 3806
rect 222292 3742 222344 3748
rect 223408 3534 223436 6052
rect 223396 3528 223448 3534
rect 223396 3470 223448 3476
rect 223948 3188 224000 3194
rect 223948 3130 224000 3136
rect 221556 3120 221608 3126
rect 221556 3062 221608 3068
rect 221188 3052 221240 3058
rect 221188 2994 221240 3000
rect 220452 2984 220504 2990
rect 220452 2926 220504 2932
rect 220464 480 220492 2926
rect 221568 480 221596 3062
rect 222752 3052 222804 3058
rect 222752 2994 222804 3000
rect 222764 480 222792 2994
rect 223960 480 223988 3130
rect 224512 2990 224540 6052
rect 225616 3126 225644 6052
rect 225604 3120 225656 3126
rect 225604 3062 225656 3068
rect 226340 3120 226392 3126
rect 226340 3062 226392 3068
rect 224500 2984 224552 2990
rect 224500 2926 224552 2932
rect 225144 2984 225196 2990
rect 225144 2926 225196 2932
rect 225156 480 225184 2926
rect 226352 480 226380 3062
rect 226720 3058 226748 6052
rect 227824 3194 227852 6052
rect 228732 3732 228784 3738
rect 228732 3674 228784 3680
rect 227812 3188 227864 3194
rect 227812 3130 227864 3136
rect 226708 3052 226760 3058
rect 226708 2994 226760 3000
rect 227536 3052 227588 3058
rect 227536 2994 227588 3000
rect 227548 480 227576 2994
rect 228744 480 228772 3674
rect 228928 2990 228956 6052
rect 229836 3188 229888 3194
rect 229836 3130 229888 3136
rect 228916 2984 228968 2990
rect 228916 2926 228968 2932
rect 229848 480 229876 3130
rect 230032 3126 230060 6052
rect 230020 3120 230072 3126
rect 230020 3062 230072 3068
rect 231032 3120 231084 3126
rect 231032 3062 231084 3068
rect 231044 480 231072 3062
rect 231136 3058 231164 6052
rect 232240 3738 232268 6052
rect 232228 3732 232280 3738
rect 232228 3674 232280 3680
rect 233344 3194 233372 6052
rect 233332 3188 233384 3194
rect 233332 3130 233384 3136
rect 234448 3126 234476 6052
rect 234436 3120 234488 3126
rect 234436 3062 234488 3068
rect 234620 3120 234672 3126
rect 234620 3062 234672 3068
rect 231124 3052 231176 3058
rect 231124 2994 231176 3000
rect 233424 3052 233476 3058
rect 233424 2994 233476 3000
rect 232228 2984 232280 2990
rect 232228 2926 232280 2932
rect 232240 480 232268 2926
rect 233436 480 233464 2994
rect 234632 480 234660 3062
rect 235552 2990 235580 6052
rect 236656 3058 236684 6052
rect 237760 3126 237788 6052
rect 237748 3120 237800 3126
rect 237748 3062 237800 3068
rect 238116 3120 238168 3126
rect 238116 3062 238168 3068
rect 236644 3052 236696 3058
rect 236644 2994 236696 3000
rect 237012 3052 237064 3058
rect 237012 2994 237064 3000
rect 235540 2984 235592 2990
rect 235540 2926 235592 2932
rect 235816 2916 235868 2922
rect 235816 2858 235868 2864
rect 235828 480 235856 2858
rect 237024 480 237052 2994
rect 238128 480 238156 3062
rect 238864 2922 238892 6052
rect 239968 3058 239996 6052
rect 241072 3126 241100 6052
rect 241060 3120 241112 3126
rect 241060 3062 241112 3068
rect 241704 3120 241756 3126
rect 241704 3062 241756 3068
rect 239956 3052 240008 3058
rect 239956 2994 240008 3000
rect 240508 3052 240560 3058
rect 240508 2994 240560 3000
rect 239312 2984 239364 2990
rect 239312 2926 239364 2932
rect 238852 2916 238904 2922
rect 238852 2858 238904 2864
rect 239324 480 239352 2926
rect 240520 480 240548 2994
rect 241716 480 241744 3062
rect 242176 2990 242204 6052
rect 243280 3058 243308 6052
rect 244384 3126 244412 6052
rect 244372 3120 244424 3126
rect 244372 3062 244424 3068
rect 243268 3052 243320 3058
rect 243268 2994 243320 3000
rect 244096 3052 244148 3058
rect 244096 2994 244148 3000
rect 242164 2984 242216 2990
rect 242164 2926 242216 2932
rect 242900 2916 242952 2922
rect 242900 2858 242952 2864
rect 242912 480 242940 2858
rect 244108 480 244136 2994
rect 245200 2984 245252 2990
rect 245200 2926 245252 2932
rect 245212 480 245240 2926
rect 245488 2922 245516 6052
rect 246396 3188 246448 3194
rect 246396 3130 246448 3136
rect 245476 2916 245528 2922
rect 245476 2858 245528 2864
rect 246408 480 246436 3130
rect 246592 3058 246620 6052
rect 247592 3120 247644 3126
rect 247592 3062 247644 3068
rect 246580 3052 246632 3058
rect 246580 2994 246632 3000
rect 247604 480 247632 3062
rect 247696 2990 247724 6052
rect 248800 3194 248828 6052
rect 248788 3188 248840 3194
rect 248788 3130 248840 3136
rect 249904 3126 249932 6052
rect 249892 3120 249944 3126
rect 249892 3062 249944 3068
rect 249984 3120 250036 3126
rect 249984 3062 250036 3068
rect 248788 3052 248840 3058
rect 248788 2994 248840 3000
rect 247684 2984 247736 2990
rect 247684 2926 247736 2932
rect 248800 480 248828 2994
rect 249996 480 250024 3062
rect 251008 3058 251036 6052
rect 252112 3126 252140 6052
rect 252100 3120 252152 3126
rect 252100 3062 252152 3068
rect 252376 3120 252428 3126
rect 252376 3062 252428 3068
rect 250996 3052 251048 3058
rect 250996 2994 251048 3000
rect 251180 3052 251232 3058
rect 251180 2994 251232 3000
rect 251192 480 251220 2994
rect 252388 480 252416 3062
rect 253216 3058 253244 6052
rect 254320 3126 254348 6052
rect 254308 3120 254360 3126
rect 254308 3062 254360 3068
rect 254676 3120 254728 3126
rect 254676 3062 254728 3068
rect 253204 3052 253256 3058
rect 253204 2994 253256 3000
rect 253480 3052 253532 3058
rect 253480 2994 253532 3000
rect 253492 480 253520 2994
rect 254688 480 254716 3062
rect 255424 3058 255452 6052
rect 256528 3126 256556 6052
rect 256516 3120 256568 3126
rect 256516 3062 256568 3068
rect 257068 3120 257120 3126
rect 257068 3062 257120 3068
rect 255412 3052 255464 3058
rect 255412 2994 255464 3000
rect 255872 3052 255924 3058
rect 255872 2994 255924 3000
rect 255884 480 255912 2994
rect 257080 480 257108 3062
rect 257632 3058 257660 6052
rect 258736 3126 258764 6052
rect 258724 3120 258776 3126
rect 258724 3062 258776 3068
rect 259460 3120 259512 3126
rect 259460 3062 259512 3068
rect 257620 3052 257672 3058
rect 257620 2994 257672 3000
rect 258264 3052 258316 3058
rect 258264 2994 258316 3000
rect 258276 480 258304 2994
rect 259472 480 259500 3062
rect 259840 3058 259868 6052
rect 260944 3126 260972 6052
rect 260932 3120 260984 3126
rect 260932 3062 260984 3068
rect 261760 3120 261812 3126
rect 261760 3062 261812 3068
rect 259828 3052 259880 3058
rect 259828 2994 259880 3000
rect 260656 3052 260708 3058
rect 260656 2994 260708 3000
rect 260668 480 260696 2994
rect 261772 480 261800 3062
rect 262048 3058 262076 6052
rect 263152 3126 263180 6052
rect 263140 3120 263192 3126
rect 263140 3062 263192 3068
rect 264152 3120 264204 3126
rect 264152 3062 264204 3068
rect 262036 3052 262088 3058
rect 262036 2994 262088 3000
rect 262956 3052 263008 3058
rect 262956 2994 263008 3000
rect 262968 480 262996 2994
rect 264164 480 264192 3062
rect 264256 3058 264284 6052
rect 265360 3126 265388 6052
rect 265348 3120 265400 3126
rect 265348 3062 265400 3068
rect 264244 3052 264296 3058
rect 264244 2994 264296 3000
rect 266464 2922 266492 6052
rect 267016 6038 267582 6066
rect 265348 2916 265400 2922
rect 265348 2858 265400 2864
rect 266452 2916 266504 2922
rect 266452 2858 266504 2864
rect 265360 480 265388 2858
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 354 266626 480
rect 267016 354 267044 6038
rect 268672 3058 268700 6052
rect 267740 3052 267792 3058
rect 267740 2994 267792 3000
rect 268660 3052 268712 3058
rect 268660 2994 268712 3000
rect 267752 480 267780 2994
rect 269776 2922 269804 6052
rect 270512 6038 270894 6066
rect 268844 2916 268896 2922
rect 268844 2858 268896 2864
rect 269764 2916 269816 2922
rect 269764 2858 269816 2864
rect 268856 480 268884 2858
rect 270512 2802 270540 6038
rect 271984 3126 272012 6052
rect 272720 6038 273102 6066
rect 273640 6038 274206 6066
rect 275020 6038 275310 6066
rect 276032 6038 276414 6066
rect 277412 6038 277518 6066
rect 278332 6038 278622 6066
rect 279528 6038 279726 6066
rect 280724 6038 280830 6066
rect 271236 3120 271288 3126
rect 271236 3062 271288 3068
rect 271972 3120 272024 3126
rect 271972 3062 272024 3068
rect 270420 2774 270540 2802
rect 266514 326 267044 354
rect 266514 -960 266626 326
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 354 270122 480
rect 270420 354 270448 2774
rect 271248 480 271276 3062
rect 270010 326 270448 354
rect 270010 -960 270122 326
rect 271206 -960 271318 480
rect 272402 354 272514 480
rect 272720 354 272748 6038
rect 273640 480 273668 6038
rect 272402 326 272748 354
rect 272402 -960 272514 326
rect 273598 -960 273710 480
rect 274794 218 274906 480
rect 275020 218 275048 6038
rect 276032 480 276060 6038
rect 277412 3074 277440 6038
rect 277136 3046 277440 3074
rect 277136 480 277164 3046
rect 278332 480 278360 6038
rect 279528 480 279556 6038
rect 280724 480 280752 6038
rect 281920 480 281948 6052
rect 283038 6038 283144 6066
rect 284142 6038 284248 6066
rect 285246 6038 285444 6066
rect 286350 6038 286640 6066
rect 283116 480 283144 6038
rect 284220 3074 284248 6038
rect 284220 3046 284340 3074
rect 284312 480 284340 3046
rect 285416 480 285444 6038
rect 286612 480 286640 6038
rect 274794 190 275048 218
rect 274794 -960 274906 190
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287440 354 287468 6052
rect 288558 6038 289032 6066
rect 289662 6038 289768 6066
rect 290766 6038 291148 6066
rect 289004 480 289032 6038
rect 289740 2802 289768 6038
rect 291120 3074 291148 6038
rect 291120 3046 291424 3074
rect 291856 3058 291884 6052
rect 292974 6038 293264 6066
rect 289740 2774 289860 2802
rect 287766 354 287878 480
rect 287440 326 287878 354
rect 287766 -960 287878 326
rect 288962 -960 289074 480
rect 289832 354 289860 2774
rect 291396 480 291424 3046
rect 291844 3052 291896 3058
rect 291844 2994 291896 3000
rect 292580 3052 292632 3058
rect 292580 2994 292632 3000
rect 292592 480 292620 2994
rect 290158 354 290270 480
rect 289832 326 290270 354
rect 290158 -960 290270 326
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293236 354 293264 6038
rect 294064 3058 294092 6052
rect 295168 3058 295196 6052
rect 296272 3058 296300 6052
rect 297376 3058 297404 6052
rect 298480 3194 298508 6052
rect 298468 3188 298520 3194
rect 298468 3130 298520 3136
rect 299584 3058 299612 6052
rect 299664 3188 299716 3194
rect 299664 3130 299716 3136
rect 294052 3052 294104 3058
rect 294052 2994 294104 3000
rect 294880 3052 294932 3058
rect 294880 2994 294932 3000
rect 295156 3052 295208 3058
rect 295156 2994 295208 3000
rect 296076 3052 296128 3058
rect 296076 2994 296128 3000
rect 296260 3052 296312 3058
rect 296260 2994 296312 3000
rect 297272 3052 297324 3058
rect 297272 2994 297324 3000
rect 297364 3052 297416 3058
rect 297364 2994 297416 3000
rect 298468 3052 298520 3058
rect 298468 2994 298520 3000
rect 299572 3052 299624 3058
rect 299572 2994 299624 3000
rect 294892 480 294920 2994
rect 296088 480 296116 2994
rect 297284 480 297312 2994
rect 298480 480 298508 2994
rect 299676 480 299704 3130
rect 300688 3126 300716 6052
rect 300676 3120 300728 3126
rect 300676 3062 300728 3068
rect 301792 3058 301820 6052
rect 302896 3126 302924 6052
rect 301964 3120 302016 3126
rect 301964 3062 302016 3068
rect 302884 3120 302936 3126
rect 302884 3062 302936 3068
rect 300768 3052 300820 3058
rect 300768 2994 300820 3000
rect 301780 3052 301832 3058
rect 301780 2994 301832 3000
rect 300780 480 300808 2994
rect 301976 480 302004 3062
rect 304000 3058 304028 6052
rect 305104 3126 305132 6052
rect 304356 3120 304408 3126
rect 304356 3062 304408 3068
rect 305092 3120 305144 3126
rect 305092 3062 305144 3068
rect 303160 3052 303212 3058
rect 303160 2994 303212 3000
rect 303988 3052 304040 3058
rect 303988 2994 304040 3000
rect 303172 480 303200 2994
rect 304368 480 304396 3062
rect 306208 3058 306236 6052
rect 307312 3126 307340 6052
rect 306748 3120 306800 3126
rect 306748 3062 306800 3068
rect 307300 3120 307352 3126
rect 307300 3062 307352 3068
rect 305552 3052 305604 3058
rect 305552 2994 305604 3000
rect 306196 3052 306248 3058
rect 306196 2994 306248 3000
rect 305564 480 305592 2994
rect 306760 480 306788 3062
rect 308416 3058 308444 6052
rect 309048 3120 309100 3126
rect 309048 3062 309100 3068
rect 307944 3052 307996 3058
rect 307944 2994 307996 3000
rect 308404 3052 308456 3058
rect 308404 2994 308456 3000
rect 307956 480 307984 2994
rect 309060 480 309088 3062
rect 309520 2854 309548 6052
rect 310624 3058 310652 6052
rect 311728 3126 311756 6052
rect 311716 3120 311768 3126
rect 311716 3062 311768 3068
rect 310244 3052 310296 3058
rect 310244 2994 310296 3000
rect 310612 3052 310664 3058
rect 310612 2994 310664 3000
rect 312636 3052 312688 3058
rect 312636 2994 312688 3000
rect 309508 2848 309560 2854
rect 309508 2790 309560 2796
rect 310256 480 310284 2994
rect 311440 2848 311492 2854
rect 311440 2790 311492 2796
rect 311452 480 311480 2790
rect 312648 480 312676 2994
rect 312832 2854 312860 6052
rect 313832 3120 313884 3126
rect 313832 3062 313884 3068
rect 312820 2848 312872 2854
rect 312820 2790 312872 2796
rect 313844 480 313872 3062
rect 313936 3058 313964 6052
rect 315040 3126 315068 6052
rect 315028 3120 315080 3126
rect 315028 3062 315080 3068
rect 313924 3052 313976 3058
rect 313924 2994 313976 3000
rect 316144 2990 316172 6052
rect 317248 3058 317276 6052
rect 317328 3120 317380 3126
rect 317328 3062 317380 3068
rect 316224 3052 316276 3058
rect 316224 2994 316276 3000
rect 317236 3052 317288 3058
rect 317236 2994 317288 3000
rect 316132 2984 316184 2990
rect 316132 2926 316184 2932
rect 315028 2848 315080 2854
rect 315028 2790 315080 2796
rect 315040 480 315068 2790
rect 316236 480 316264 2994
rect 317340 480 317368 3062
rect 318352 2854 318380 6052
rect 319456 3126 319484 6052
rect 319444 3120 319496 3126
rect 319444 3062 319496 3068
rect 320560 3058 320588 6052
rect 319720 3052 319772 3058
rect 319720 2994 319772 3000
rect 320548 3052 320600 3058
rect 320548 2994 320600 3000
rect 318524 2984 318576 2990
rect 318524 2926 318576 2932
rect 318340 2848 318392 2854
rect 318340 2790 318392 2796
rect 318536 480 318564 2926
rect 319732 480 319760 2994
rect 321664 2854 321692 6052
rect 322768 3194 322796 6052
rect 322756 3188 322808 3194
rect 322756 3130 322808 3136
rect 322112 3120 322164 3126
rect 322112 3062 322164 3068
rect 320916 2848 320968 2854
rect 320916 2790 320968 2796
rect 321652 2848 321704 2854
rect 321652 2790 321704 2796
rect 320928 480 320956 2790
rect 322124 480 322152 3062
rect 323308 3052 323360 3058
rect 323308 2994 323360 3000
rect 323320 480 323348 2994
rect 323872 2990 323900 6052
rect 324976 3126 325004 6052
rect 325608 3188 325660 3194
rect 325608 3130 325660 3136
rect 324964 3120 325016 3126
rect 324964 3062 325016 3068
rect 323860 2984 323912 2990
rect 323860 2926 323912 2932
rect 324412 2848 324464 2854
rect 324412 2790 324464 2796
rect 324424 480 324452 2790
rect 325620 480 325648 3130
rect 326080 3058 326108 6052
rect 326068 3052 326120 3058
rect 326068 2994 326120 3000
rect 327184 2990 327212 6052
rect 328288 3126 328316 6052
rect 328000 3120 328052 3126
rect 328000 3062 328052 3068
rect 328276 3120 328328 3126
rect 328276 3062 328328 3068
rect 326804 2984 326856 2990
rect 326804 2926 326856 2932
rect 327172 2984 327224 2990
rect 327172 2926 327224 2932
rect 326816 480 326844 2926
rect 328012 480 328040 3062
rect 329196 3052 329248 3058
rect 329196 2994 329248 3000
rect 329208 480 329236 2994
rect 329392 2922 329420 6052
rect 330496 3058 330524 6052
rect 331600 3262 331628 6052
rect 331588 3256 331640 3262
rect 331588 3198 331640 3204
rect 332704 3126 332732 6052
rect 331588 3120 331640 3126
rect 331588 3062 331640 3068
rect 332692 3120 332744 3126
rect 332692 3062 332744 3068
rect 330484 3052 330536 3058
rect 330484 2994 330536 3000
rect 330392 2984 330444 2990
rect 330392 2926 330444 2932
rect 329380 2916 329432 2922
rect 329380 2858 329432 2864
rect 330404 480 330432 2926
rect 331600 480 331628 3062
rect 333808 2990 333836 6052
rect 334912 3602 334940 6052
rect 334900 3596 334952 3602
rect 334900 3538 334952 3544
rect 335084 3256 335136 3262
rect 335084 3198 335136 3204
rect 333888 3052 333940 3058
rect 333888 2994 333940 3000
rect 333796 2984 333848 2990
rect 333796 2926 333848 2932
rect 332692 2916 332744 2922
rect 332692 2858 332744 2864
rect 332704 480 332732 2858
rect 333900 480 333928 2994
rect 335096 480 335124 3198
rect 336016 3058 336044 6052
rect 337120 3126 337148 6052
rect 336280 3120 336332 3126
rect 336280 3062 336332 3068
rect 337108 3120 337160 3126
rect 337108 3062 337160 3068
rect 336004 3052 336056 3058
rect 336004 2994 336056 3000
rect 336292 480 336320 3062
rect 338224 2990 338252 6052
rect 338672 3596 338724 3602
rect 338672 3538 338724 3544
rect 337476 2984 337528 2990
rect 337476 2926 337528 2932
rect 338212 2984 338264 2990
rect 338212 2926 338264 2932
rect 337488 480 337516 2926
rect 338684 480 338712 3538
rect 339328 2922 339356 6052
rect 340432 3058 340460 6052
rect 341536 3194 341564 6052
rect 341524 3188 341576 3194
rect 341524 3130 341576 3136
rect 340972 3120 341024 3126
rect 340972 3062 341024 3068
rect 339868 3052 339920 3058
rect 339868 2994 339920 3000
rect 340420 3052 340472 3058
rect 340420 2994 340472 3000
rect 339316 2916 339368 2922
rect 339316 2858 339368 2864
rect 339880 480 339908 2994
rect 340984 480 341012 3062
rect 342640 2990 342668 6052
rect 343744 3670 343772 6052
rect 343732 3664 343784 3670
rect 343732 3606 343784 3612
rect 344848 3466 344876 6052
rect 344836 3460 344888 3466
rect 344836 3402 344888 3408
rect 345756 3188 345808 3194
rect 345756 3130 345808 3136
rect 344560 3052 344612 3058
rect 344560 2994 344612 3000
rect 342168 2984 342220 2990
rect 342168 2926 342220 2932
rect 342628 2984 342680 2990
rect 342628 2926 342680 2932
rect 342180 480 342208 2926
rect 343364 2916 343416 2922
rect 343364 2858 343416 2864
rect 343376 480 343404 2858
rect 344572 480 344600 2994
rect 345768 480 345796 3130
rect 345952 3126 345980 6052
rect 345940 3120 345992 3126
rect 345940 3062 345992 3068
rect 347056 3058 347084 6052
rect 348056 3664 348108 3670
rect 348056 3606 348108 3612
rect 347044 3052 347096 3058
rect 347044 2994 347096 3000
rect 346952 2984 347004 2990
rect 346952 2926 347004 2932
rect 346964 480 346992 2926
rect 348068 480 348096 3606
rect 348160 3194 348188 6052
rect 349264 3602 349292 6052
rect 349252 3596 349304 3602
rect 349252 3538 349304 3544
rect 349252 3460 349304 3466
rect 349252 3402 349304 3408
rect 348148 3188 348200 3194
rect 348148 3130 348200 3136
rect 349264 480 349292 3402
rect 350368 2922 350396 6052
rect 350448 3120 350500 3126
rect 350448 3062 350500 3068
rect 350356 2916 350408 2922
rect 350356 2858 350408 2864
rect 350460 480 350488 3062
rect 351472 2990 351500 6052
rect 352576 3466 352604 6052
rect 353680 3874 353708 6052
rect 353668 3868 353720 3874
rect 353668 3810 353720 3816
rect 354036 3596 354088 3602
rect 354036 3538 354088 3544
rect 352564 3460 352616 3466
rect 352564 3402 352616 3408
rect 352840 3188 352892 3194
rect 352840 3130 352892 3136
rect 351644 3052 351696 3058
rect 351644 2994 351696 3000
rect 351460 2984 351512 2990
rect 351460 2926 351512 2932
rect 351656 480 351684 2994
rect 352852 480 352880 3130
rect 354048 480 354076 3538
rect 354784 3058 354812 6052
rect 354772 3052 354824 3058
rect 354772 2994 354824 3000
rect 355888 2922 355916 6052
rect 356992 3262 357020 6052
rect 357532 3460 357584 3466
rect 357532 3402 357584 3408
rect 356980 3256 357032 3262
rect 356980 3198 357032 3204
rect 356336 2984 356388 2990
rect 356336 2926 356388 2932
rect 355232 2916 355284 2922
rect 355232 2858 355284 2864
rect 355876 2916 355928 2922
rect 355876 2858 355928 2864
rect 355244 480 355272 2858
rect 356348 480 356376 2926
rect 357544 480 357572 3402
rect 358096 2854 358124 6052
rect 358728 3868 358780 3874
rect 358728 3810 358780 3816
rect 358084 2848 358136 2854
rect 358084 2790 358136 2796
rect 358740 480 358768 3810
rect 359200 3126 359228 6052
rect 360304 3194 360332 6052
rect 360292 3188 360344 3194
rect 360292 3130 360344 3136
rect 359188 3120 359240 3126
rect 359188 3062 359240 3068
rect 359924 3052 359976 3058
rect 359924 2994 359976 3000
rect 359936 480 359964 2994
rect 361408 2990 361436 6052
rect 362512 3466 362540 6052
rect 363616 3670 363644 6052
rect 363604 3664 363656 3670
rect 363604 3606 363656 3612
rect 362500 3460 362552 3466
rect 362500 3402 362552 3408
rect 362316 3256 362368 3262
rect 362316 3198 362368 3204
rect 361396 2984 361448 2990
rect 361396 2926 361448 2932
rect 361120 2916 361172 2922
rect 361120 2858 361172 2864
rect 361132 480 361160 2858
rect 362328 480 362356 3198
rect 364616 3120 364668 3126
rect 364616 3062 364668 3068
rect 363512 2848 363564 2854
rect 363512 2790 363564 2796
rect 363524 480 363552 2790
rect 364628 480 364656 3062
rect 364720 3058 364748 6052
rect 365824 3330 365852 6052
rect 365812 3324 365864 3330
rect 365812 3266 365864 3272
rect 365812 3188 365864 3194
rect 365812 3130 365864 3136
rect 364708 3052 364760 3058
rect 364708 2994 364760 3000
rect 365824 480 365852 3130
rect 366928 2854 366956 6052
rect 368032 2990 368060 6052
rect 368204 3460 368256 3466
rect 368204 3402 368256 3408
rect 367008 2984 367060 2990
rect 367008 2926 367060 2932
rect 368020 2984 368072 2990
rect 368020 2926 368072 2932
rect 366916 2848 366968 2854
rect 366916 2790 366968 2796
rect 367020 480 367048 2926
rect 368216 480 368244 3402
rect 369136 3126 369164 6052
rect 369400 3664 369452 3670
rect 369400 3606 369452 3612
rect 369124 3120 369176 3126
rect 369124 3062 369176 3068
rect 369412 480 369440 3606
rect 370240 3194 370268 6052
rect 371344 3874 371372 6052
rect 371332 3868 371384 3874
rect 371332 3810 371384 3816
rect 372448 3534 372476 6052
rect 373552 3602 373580 6052
rect 373540 3596 373592 3602
rect 373540 3538 373592 3544
rect 372436 3528 372488 3534
rect 372436 3470 372488 3476
rect 371700 3324 371752 3330
rect 371700 3266 371752 3272
rect 370228 3188 370280 3194
rect 370228 3130 370280 3136
rect 370596 3052 370648 3058
rect 370596 2994 370648 3000
rect 370608 480 370636 2994
rect 371712 480 371740 3266
rect 374656 3058 374684 6052
rect 375288 3120 375340 3126
rect 375288 3062 375340 3068
rect 374644 3052 374696 3058
rect 374644 2994 374696 3000
rect 374092 2984 374144 2990
rect 374092 2926 374144 2932
rect 372896 2848 372948 2854
rect 372896 2790 372948 2796
rect 372908 480 372936 2790
rect 374104 480 374132 2926
rect 375300 480 375328 3062
rect 375760 2922 375788 6052
rect 376864 3194 376892 6052
rect 377680 3868 377732 3874
rect 377680 3810 377732 3816
rect 376484 3188 376536 3194
rect 376484 3130 376536 3136
rect 376852 3188 376904 3194
rect 376852 3130 376904 3136
rect 375748 2916 375800 2922
rect 375748 2858 375800 2864
rect 376496 480 376524 3130
rect 377692 480 377720 3810
rect 377968 2990 377996 6052
rect 378876 3528 378928 3534
rect 378876 3470 378928 3476
rect 377956 2984 378008 2990
rect 377956 2926 378008 2932
rect 378888 480 378916 3470
rect 379072 3126 379100 6052
rect 380176 3670 380204 6052
rect 381280 3806 381308 6052
rect 381268 3800 381320 3806
rect 381268 3742 381320 3748
rect 380164 3664 380216 3670
rect 380164 3606 380216 3612
rect 382384 3602 382412 6052
rect 379980 3596 380032 3602
rect 379980 3538 380032 3544
rect 382372 3596 382424 3602
rect 382372 3538 382424 3544
rect 379060 3120 379112 3126
rect 379060 3062 379112 3068
rect 379992 480 380020 3538
rect 383488 3466 383516 6052
rect 383476 3460 383528 3466
rect 383476 3402 383528 3408
rect 384592 3194 384620 6052
rect 383568 3188 383620 3194
rect 383568 3130 383620 3136
rect 384580 3188 384632 3194
rect 384580 3130 384632 3136
rect 381176 3052 381228 3058
rect 381176 2994 381228 3000
rect 381188 480 381216 2994
rect 382372 2916 382424 2922
rect 382372 2858 382424 2864
rect 382384 480 382412 2858
rect 383580 480 383608 3130
rect 385696 2990 385724 6052
rect 386800 3126 386828 6052
rect 387156 3664 387208 3670
rect 387156 3606 387208 3612
rect 385960 3120 386012 3126
rect 385960 3062 386012 3068
rect 386788 3120 386840 3126
rect 386788 3062 386840 3068
rect 384764 2984 384816 2990
rect 384764 2926 384816 2932
rect 385684 2984 385736 2990
rect 385684 2926 385736 2932
rect 384776 480 384804 2926
rect 385972 480 386000 3062
rect 387168 480 387196 3606
rect 387904 3058 387932 6052
rect 388260 3800 388312 3806
rect 388260 3742 388312 3748
rect 387892 3052 387944 3058
rect 387892 2994 387944 3000
rect 388272 480 388300 3742
rect 389008 3534 389036 6052
rect 390112 3602 390140 6052
rect 391216 3670 391244 6052
rect 391204 3664 391256 3670
rect 391204 3606 391256 3612
rect 389456 3596 389508 3602
rect 389456 3538 389508 3544
rect 390100 3596 390152 3602
rect 390100 3538 390152 3544
rect 388996 3528 389048 3534
rect 388996 3470 389048 3476
rect 389468 480 389496 3538
rect 390652 3460 390704 3466
rect 390652 3402 390704 3408
rect 390664 480 390692 3402
rect 392320 3398 392348 6052
rect 392308 3392 392360 3398
rect 392308 3334 392360 3340
rect 393424 3194 393452 6052
rect 391848 3188 391900 3194
rect 391848 3130 391900 3136
rect 393412 3188 393464 3194
rect 393412 3130 393464 3136
rect 391860 480 391888 3130
rect 394240 3120 394292 3126
rect 394240 3062 394292 3068
rect 393044 2984 393096 2990
rect 393044 2926 393096 2932
rect 393056 480 393084 2926
rect 394252 480 394280 3062
rect 394528 2990 394556 6052
rect 395632 3466 395660 6052
rect 396540 3528 396592 3534
rect 396540 3470 396592 3476
rect 395620 3460 395672 3466
rect 395620 3402 395672 3408
rect 395344 3052 395396 3058
rect 395344 2994 395396 3000
rect 394516 2984 394568 2990
rect 394516 2926 394568 2932
rect 395356 480 395384 2994
rect 396552 480 396580 3470
rect 396736 3058 396764 6052
rect 397840 3874 397868 6052
rect 397828 3868 397880 3874
rect 397828 3810 397880 3816
rect 398944 3806 398972 6052
rect 400048 4078 400076 6052
rect 400036 4072 400088 4078
rect 400036 4014 400088 4020
rect 401152 3942 401180 6052
rect 401140 3936 401192 3942
rect 401140 3878 401192 3884
rect 398932 3800 398984 3806
rect 398932 3742 398984 3748
rect 398932 3664 398984 3670
rect 398932 3606 398984 3612
rect 397736 3596 397788 3602
rect 397736 3538 397788 3544
rect 396724 3052 396776 3058
rect 396724 2994 396776 3000
rect 397748 480 397776 3538
rect 398944 480 398972 3606
rect 402256 3602 402284 6052
rect 402244 3596 402296 3602
rect 402244 3538 402296 3544
rect 400128 3392 400180 3398
rect 400128 3334 400180 3340
rect 400140 480 400168 3334
rect 401324 3188 401376 3194
rect 401324 3130 401376 3136
rect 401336 480 401364 3130
rect 403360 3126 403388 6052
rect 404464 3534 404492 6052
rect 405568 3670 405596 6052
rect 406016 3868 406068 3874
rect 406016 3810 406068 3816
rect 405556 3664 405608 3670
rect 405556 3606 405608 3612
rect 404452 3528 404504 3534
rect 404452 3470 404504 3476
rect 403624 3460 403676 3466
rect 403624 3402 403676 3408
rect 403348 3120 403400 3126
rect 403348 3062 403400 3068
rect 402520 2984 402572 2990
rect 402520 2926 402572 2932
rect 402532 480 402560 2926
rect 403636 480 403664 3402
rect 404820 3052 404872 3058
rect 404820 2994 404872 3000
rect 404832 480 404860 2994
rect 406028 480 406056 3810
rect 406672 3466 406700 6052
rect 407776 4010 407804 6052
rect 408408 4072 408460 4078
rect 408408 4014 408460 4020
rect 407764 4004 407816 4010
rect 407764 3946 407816 3952
rect 407212 3800 407264 3806
rect 407212 3742 407264 3748
rect 406660 3460 406712 3466
rect 406660 3402 406712 3408
rect 407224 480 407252 3742
rect 408420 480 408448 4014
rect 408880 3942 408908 6052
rect 408868 3936 408920 3942
rect 408868 3878 408920 3884
rect 409984 3874 410012 6052
rect 409604 3868 409656 3874
rect 409604 3810 409656 3816
rect 409972 3868 410024 3874
rect 409972 3810 410024 3816
rect 409616 480 409644 3810
rect 411088 3806 411116 6052
rect 411076 3800 411128 3806
rect 411076 3742 411128 3748
rect 412192 3602 412220 6052
rect 410800 3596 410852 3602
rect 410800 3538 410852 3544
rect 412180 3596 412232 3602
rect 412180 3538 412232 3544
rect 410812 480 410840 3538
rect 413100 3528 413152 3534
rect 413100 3470 413152 3476
rect 411904 3120 411956 3126
rect 411904 3062 411956 3068
rect 411916 480 411944 3062
rect 413112 480 413140 3470
rect 413296 3398 413324 6052
rect 414400 3670 414428 6052
rect 415504 4146 415532 6052
rect 415492 4140 415544 4146
rect 415492 4082 415544 4088
rect 416608 4010 416636 6052
rect 416596 4004 416648 4010
rect 416596 3946 416648 3952
rect 417712 3942 417740 6052
rect 416688 3936 416740 3942
rect 416688 3878 416740 3884
rect 417700 3936 417752 3942
rect 417700 3878 417752 3884
rect 414296 3664 414348 3670
rect 414296 3606 414348 3612
rect 414388 3664 414440 3670
rect 414388 3606 414440 3612
rect 413284 3392 413336 3398
rect 413284 3334 413336 3340
rect 414308 480 414336 3606
rect 415492 3460 415544 3466
rect 415492 3402 415544 3408
rect 415504 480 415532 3402
rect 416700 480 416728 3878
rect 417884 3868 417936 3874
rect 417884 3810 417936 3816
rect 417896 480 417924 3810
rect 418816 3330 418844 6052
rect 418988 3800 419040 3806
rect 418988 3742 419040 3748
rect 418804 3324 418856 3330
rect 418804 3266 418856 3272
rect 419000 480 419028 3742
rect 419920 3534 419948 6052
rect 421024 4078 421052 6052
rect 421012 4072 421064 4078
rect 421012 4014 421064 4020
rect 420184 3732 420236 3738
rect 420184 3674 420236 3680
rect 419908 3528 419960 3534
rect 419908 3470 419960 3476
rect 420196 480 420224 3674
rect 422128 3602 422156 6052
rect 423232 3806 423260 6052
rect 424336 3874 424364 6052
rect 424968 4140 425020 4146
rect 424968 4082 425020 4088
rect 424324 3868 424376 3874
rect 424324 3810 424376 3816
rect 423220 3800 423272 3806
rect 423220 3742 423272 3748
rect 423772 3732 423824 3738
rect 423772 3674 423824 3680
rect 421380 3596 421432 3602
rect 421380 3538 421432 3544
rect 422116 3596 422168 3602
rect 422116 3538 422168 3544
rect 421392 480 421420 3538
rect 422576 3528 422628 3534
rect 422576 3470 422628 3476
rect 422588 480 422616 3470
rect 423784 480 423812 3674
rect 424980 480 425008 4082
rect 425440 3738 425468 6052
rect 426544 4010 426572 6052
rect 426164 4004 426216 4010
rect 426164 3946 426216 3952
rect 426532 4004 426584 4010
rect 426532 3946 426584 3952
rect 425428 3732 425480 3738
rect 425428 3674 425480 3680
rect 426176 480 426204 3946
rect 427648 3942 427676 6052
rect 427268 3936 427320 3942
rect 427268 3878 427320 3884
rect 427636 3936 427688 3942
rect 427636 3878 427688 3884
rect 427280 480 427308 3878
rect 428752 3534 428780 6052
rect 429660 3664 429712 3670
rect 429660 3606 429712 3612
rect 428740 3528 428792 3534
rect 428740 3470 428792 3476
rect 428464 3460 428516 3466
rect 428464 3402 428516 3408
rect 428476 480 428504 3402
rect 429672 480 429700 3606
rect 429856 3466 429884 6052
rect 430960 4146 430988 6052
rect 430948 4140 431000 4146
rect 430948 4082 431000 4088
rect 432064 4078 432092 6052
rect 430856 4072 430908 4078
rect 430856 4014 430908 4020
rect 432052 4072 432104 4078
rect 432052 4014 432104 4020
rect 429844 3460 429896 3466
rect 429844 3402 429896 3408
rect 430868 480 430896 4014
rect 433168 3602 433196 6052
rect 434286 6038 434576 6066
rect 434548 3874 434576 6038
rect 434444 3868 434496 3874
rect 434444 3810 434496 3816
rect 434536 3868 434588 3874
rect 434536 3810 434588 3816
rect 433248 3800 433300 3806
rect 433248 3742 433300 3748
rect 432052 3596 432104 3602
rect 432052 3538 432104 3544
rect 433156 3596 433208 3602
rect 433156 3538 433208 3544
rect 432064 480 432092 3538
rect 433260 480 433288 3742
rect 434456 480 434484 3810
rect 435376 3806 435404 6052
rect 435364 3800 435416 3806
rect 435364 3742 435416 3748
rect 436480 3738 436508 6052
rect 437584 4010 437612 6052
rect 436744 4004 436796 4010
rect 436744 3946 436796 3952
rect 437572 4004 437624 4010
rect 437572 3946 437624 3952
rect 435548 3732 435600 3738
rect 435548 3674 435600 3680
rect 436468 3732 436520 3738
rect 436468 3674 436520 3680
rect 435560 480 435588 3674
rect 436756 480 436784 3946
rect 437940 3936 437992 3942
rect 437940 3878 437992 3884
rect 437952 480 437980 3878
rect 438688 3398 438716 6052
rect 439792 3534 439820 6052
rect 439136 3528 439188 3534
rect 439136 3470 439188 3476
rect 439780 3528 439832 3534
rect 439780 3470 439832 3476
rect 438676 3392 438728 3398
rect 438676 3334 438728 3340
rect 439148 480 439176 3470
rect 440332 3460 440384 3466
rect 440332 3402 440384 3408
rect 440344 480 440372 3402
rect 440896 3262 440924 6052
rect 441528 4140 441580 4146
rect 441528 4082 441580 4088
rect 440884 3256 440936 3262
rect 440884 3198 440936 3204
rect 441540 480 441568 4082
rect 442000 3942 442028 6052
rect 442632 4072 442684 4078
rect 442632 4014 442684 4020
rect 441988 3936 442040 3942
rect 441988 3878 442040 3884
rect 442644 480 442672 4014
rect 443104 3670 443132 6052
rect 443092 3664 443144 3670
rect 443092 3606 443144 3612
rect 444208 3602 444236 6052
rect 445024 3868 445076 3874
rect 445024 3810 445076 3816
rect 443828 3596 443880 3602
rect 443828 3538 443880 3544
rect 444196 3596 444248 3602
rect 444196 3538 444248 3544
rect 443840 480 443868 3538
rect 445036 480 445064 3810
rect 445312 3466 445340 6052
rect 446416 3874 446444 6052
rect 446404 3868 446456 3874
rect 446404 3810 446456 3816
rect 446220 3800 446272 3806
rect 446220 3742 446272 3748
rect 445300 3460 445352 3466
rect 445300 3402 445352 3408
rect 446232 480 446260 3742
rect 447416 3732 447468 3738
rect 447416 3674 447468 3680
rect 447428 480 447456 3674
rect 447520 3330 447548 6052
rect 448624 4078 448652 6052
rect 448612 4072 448664 4078
rect 448612 4014 448664 4020
rect 448520 4004 448572 4010
rect 448520 3946 448572 3952
rect 447508 3324 447560 3330
rect 447508 3266 447560 3272
rect 448532 1986 448560 3946
rect 449728 3194 449756 6052
rect 450832 3738 450860 6052
rect 451936 3806 451964 6052
rect 451924 3800 451976 3806
rect 451924 3742 451976 3748
rect 450820 3732 450872 3738
rect 450820 3674 450872 3680
rect 453040 3534 453068 6052
rect 453304 3936 453356 3942
rect 453304 3878 453356 3884
rect 450912 3528 450964 3534
rect 450912 3470 450964 3476
rect 453028 3528 453080 3534
rect 453028 3470 453080 3476
rect 449808 3392 449860 3398
rect 449808 3334 449860 3340
rect 449716 3188 449768 3194
rect 449716 3130 449768 3136
rect 448532 1958 448652 1986
rect 448624 480 448652 1958
rect 449820 480 449848 3334
rect 450924 480 450952 3470
rect 452108 3256 452160 3262
rect 452108 3198 452160 3204
rect 452120 480 452148 3198
rect 453316 480 453344 3878
rect 454144 3262 454172 6052
rect 454500 3664 454552 3670
rect 454500 3606 454552 3612
rect 454132 3256 454184 3262
rect 454132 3198 454184 3204
rect 454512 480 454540 3606
rect 455248 3398 455276 6052
rect 456352 3670 456380 6052
rect 457456 3942 457484 6052
rect 457444 3936 457496 3942
rect 457444 3878 457496 3884
rect 458560 3874 458588 6052
rect 458088 3868 458140 3874
rect 458088 3810 458140 3816
rect 458548 3868 458600 3874
rect 458548 3810 458600 3816
rect 456340 3664 456392 3670
rect 456340 3606 456392 3612
rect 455696 3596 455748 3602
rect 455696 3538 455748 3544
rect 455236 3392 455288 3398
rect 455236 3334 455288 3340
rect 455708 480 455736 3538
rect 456892 3460 456944 3466
rect 456892 3402 456944 3408
rect 456904 480 456932 3402
rect 458100 480 458128 3810
rect 459664 3466 459692 6052
rect 460388 4072 460440 4078
rect 460388 4014 460440 4020
rect 459652 3460 459704 3466
rect 459652 3402 459704 3408
rect 459192 3324 459244 3330
rect 459192 3266 459244 3272
rect 459204 480 459232 3266
rect 460400 480 460428 4014
rect 460768 3534 460796 6052
rect 461872 4010 461900 6052
rect 461860 4004 461912 4010
rect 461860 3946 461912 3952
rect 462976 3738 463004 6052
rect 464080 4146 464108 6052
rect 464068 4140 464120 4146
rect 464068 4082 464120 4088
rect 465184 4078 465212 6052
rect 465172 4072 465224 4078
rect 465172 4014 465224 4020
rect 463976 3800 464028 3806
rect 463976 3742 464028 3748
rect 462780 3732 462832 3738
rect 462780 3674 462832 3680
rect 462964 3732 463016 3738
rect 462964 3674 463016 3680
rect 460756 3528 460808 3534
rect 460756 3470 460808 3476
rect 461584 3188 461636 3194
rect 461584 3130 461636 3136
rect 461596 480 461624 3130
rect 462792 480 462820 3674
rect 463988 480 464016 3742
rect 466288 3602 466316 6052
rect 467392 3806 467420 6052
rect 467380 3800 467432 3806
rect 467380 3742 467432 3748
rect 468496 3670 468524 6052
rect 468300 3664 468352 3670
rect 468300 3606 468352 3612
rect 468484 3664 468536 3670
rect 468484 3606 468536 3612
rect 465172 3596 465224 3602
rect 465172 3538 465224 3544
rect 466276 3596 466328 3602
rect 466276 3538 466328 3544
rect 465184 480 465212 3538
rect 467472 3392 467524 3398
rect 467472 3334 467524 3340
rect 466276 3256 466328 3262
rect 466276 3198 466328 3204
rect 466288 480 466316 3198
rect 467484 480 467512 3334
rect 293654 354 293766 480
rect 293236 326 293766 354
rect 293654 -960 293766 326
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468312 354 468340 3606
rect 469600 3398 469628 6052
rect 469864 3936 469916 3942
rect 469864 3878 469916 3884
rect 469588 3392 469640 3398
rect 469588 3334 469640 3340
rect 469876 480 469904 3878
rect 470704 3126 470732 6052
rect 471808 3942 471836 6052
rect 471796 3936 471848 3942
rect 471796 3878 471848 3884
rect 471060 3868 471112 3874
rect 471060 3810 471112 3816
rect 470692 3120 470744 3126
rect 470692 3062 470744 3068
rect 471072 480 471100 3810
rect 472256 3460 472308 3466
rect 472256 3402 472308 3408
rect 472268 480 472296 3402
rect 472912 3330 472940 6052
rect 474016 3874 474044 6052
rect 475134 6038 475516 6066
rect 474556 4004 474608 4010
rect 474556 3946 474608 3952
rect 474004 3868 474056 3874
rect 474004 3810 474056 3816
rect 473452 3528 473504 3534
rect 473452 3470 473504 3476
rect 472900 3324 472952 3330
rect 472900 3266 472952 3272
rect 473464 480 473492 3470
rect 474568 480 474596 3946
rect 475384 3800 475436 3806
rect 475384 3742 475436 3748
rect 474740 3732 474792 3738
rect 474740 3674 474792 3680
rect 474752 2854 474780 3674
rect 475396 3534 475424 3742
rect 475488 3738 475516 6038
rect 476224 4078 476252 6052
rect 477328 4146 477356 6052
rect 476948 4140 477000 4146
rect 476948 4082 477000 4088
rect 477316 4140 477368 4146
rect 477316 4082 477368 4088
rect 476212 4072 476264 4078
rect 476212 4014 476264 4020
rect 475476 3732 475528 3738
rect 475476 3674 475528 3680
rect 475384 3528 475436 3534
rect 475384 3470 475436 3476
rect 474740 2848 474792 2854
rect 474740 2790 474792 2796
rect 475752 2848 475804 2854
rect 475752 2790 475804 2796
rect 475764 480 475792 2790
rect 476960 480 476988 4082
rect 478432 4010 478460 6052
rect 478144 4004 478196 4010
rect 478144 3946 478196 3952
rect 478420 4004 478472 4010
rect 478420 3946 478472 3952
rect 478156 480 478184 3946
rect 479536 3602 479564 6052
rect 479524 3596 479576 3602
rect 479524 3538 479576 3544
rect 480536 3528 480588 3534
rect 480536 3470 480588 3476
rect 479340 3460 479392 3466
rect 479340 3402 479392 3408
rect 479352 480 479380 3402
rect 480548 480 480576 3470
rect 480640 3126 480668 6052
rect 481744 4078 481772 6052
rect 481640 4072 481692 4078
rect 481640 4014 481692 4020
rect 481732 4072 481784 4078
rect 481732 4014 481784 4020
rect 481652 3534 481680 4014
rect 482848 3806 482876 6052
rect 482836 3800 482888 3806
rect 482836 3742 482888 3748
rect 483952 3670 483980 6052
rect 481732 3664 481784 3670
rect 481732 3606 481784 3612
rect 483940 3664 483992 3670
rect 483940 3606 483992 3612
rect 481640 3528 481692 3534
rect 481640 3470 481692 3476
rect 480628 3120 480680 3126
rect 480628 3062 480680 3068
rect 481744 480 481772 3606
rect 482836 3392 482888 3398
rect 482836 3334 482888 3340
rect 482848 480 482876 3334
rect 484032 3324 484084 3330
rect 484032 3266 484084 3272
rect 484044 480 484072 3266
rect 485056 3194 485084 6052
rect 485228 3936 485280 3942
rect 485228 3878 485280 3884
rect 485044 3188 485096 3194
rect 485044 3130 485096 3136
rect 485240 480 485268 3878
rect 486160 3398 486188 6052
rect 486424 3460 486476 3466
rect 486424 3402 486476 3408
rect 486148 3392 486200 3398
rect 486148 3334 486200 3340
rect 486436 480 486464 3402
rect 487264 3330 487292 6052
rect 488368 3942 488396 6052
rect 488356 3936 488408 3942
rect 488356 3878 488408 3884
rect 487620 3868 487672 3874
rect 487620 3810 487672 3816
rect 487252 3324 487304 3330
rect 487252 3266 487304 3272
rect 487632 480 487660 3810
rect 488816 3732 488868 3738
rect 488816 3674 488868 3680
rect 488828 480 488856 3674
rect 489472 3466 489500 6052
rect 490576 3534 490604 6052
rect 491116 4140 491168 4146
rect 491116 4082 491168 4088
rect 489920 3528 489972 3534
rect 489920 3470 489972 3476
rect 490564 3528 490616 3534
rect 490564 3470 490616 3476
rect 489460 3460 489512 3466
rect 489460 3402 489512 3408
rect 489932 480 489960 3470
rect 491128 480 491156 4082
rect 491680 3806 491708 6052
rect 492312 4004 492364 4010
rect 492312 3946 492364 3952
rect 491668 3800 491720 3806
rect 491668 3742 491720 3748
rect 492324 480 492352 3946
rect 492784 3262 492812 6052
rect 493888 4146 493916 6052
rect 493876 4140 493928 4146
rect 493876 4082 493928 4088
rect 494992 3738 495020 6052
rect 495900 4072 495952 4078
rect 495900 4014 495952 4020
rect 494980 3732 495032 3738
rect 494980 3674 495032 3680
rect 493508 3596 493560 3602
rect 493508 3538 493560 3544
rect 492772 3256 492824 3262
rect 492772 3198 492824 3204
rect 493520 480 493548 3538
rect 494704 3120 494756 3126
rect 494704 3062 494756 3068
rect 494716 480 494744 3062
rect 495912 480 495940 4014
rect 496096 3602 496124 6052
rect 497200 4010 497228 6052
rect 498304 4078 498332 6052
rect 498292 4072 498344 4078
rect 498292 4014 498344 4020
rect 497188 4004 497240 4010
rect 497188 3946 497240 3952
rect 497096 3868 497148 3874
rect 497096 3810 497148 3816
rect 496084 3596 496136 3602
rect 496084 3538 496136 3544
rect 497108 480 497136 3810
rect 499408 3670 499436 6052
rect 500526 6038 500816 6066
rect 501630 6038 501920 6066
rect 498200 3664 498252 3670
rect 498200 3606 498252 3612
rect 499396 3664 499448 3670
rect 499396 3606 499448 3612
rect 498212 480 498240 3606
rect 500788 3398 500816 6038
rect 500592 3392 500644 3398
rect 500592 3334 500644 3340
rect 500776 3392 500828 3398
rect 500776 3334 500828 3340
rect 499396 3188 499448 3194
rect 499396 3130 499448 3136
rect 499408 480 499436 3130
rect 500604 480 500632 3334
rect 501892 3330 501920 6038
rect 502720 3942 502748 6052
rect 502708 3936 502760 3942
rect 502708 3878 502760 3884
rect 502984 3868 503036 3874
rect 502984 3810 503036 3816
rect 501788 3324 501840 3330
rect 501788 3266 501840 3272
rect 501880 3324 501932 3330
rect 501880 3266 501932 3272
rect 501800 480 501828 3266
rect 502996 480 503024 3810
rect 503824 3126 503852 6052
rect 504928 3806 504956 6052
rect 504916 3800 504968 3806
rect 504916 3742 504968 3748
rect 505376 3528 505428 3534
rect 505376 3470 505428 3476
rect 504180 3460 504232 3466
rect 504180 3402 504232 3408
rect 503812 3120 503864 3126
rect 503812 3062 503864 3068
rect 504192 480 504220 3402
rect 505388 480 505416 3470
rect 506032 3466 506060 6052
rect 506480 3868 506532 3874
rect 506480 3810 506532 3816
rect 506020 3460 506072 3466
rect 506020 3402 506072 3408
rect 506492 480 506520 3810
rect 507136 3534 507164 6052
rect 507124 3528 507176 3534
rect 507124 3470 507176 3476
rect 507676 3256 507728 3262
rect 507676 3198 507728 3204
rect 507688 480 507716 3198
rect 508240 3058 508268 6052
rect 508872 4140 508924 4146
rect 508872 4082 508924 4088
rect 508228 3052 508280 3058
rect 508228 2994 508280 3000
rect 508884 480 508912 4082
rect 509344 3262 509372 6052
rect 510448 4146 510476 6052
rect 510436 4140 510488 4146
rect 510436 4082 510488 4088
rect 511552 3738 511580 6052
rect 512460 4004 512512 4010
rect 512460 3946 512512 3952
rect 510068 3732 510120 3738
rect 510068 3674 510120 3680
rect 511540 3732 511592 3738
rect 511540 3674 511592 3680
rect 509332 3256 509384 3262
rect 509332 3198 509384 3204
rect 510080 480 510108 3674
rect 511264 3596 511316 3602
rect 511264 3538 511316 3544
rect 511276 480 511304 3538
rect 512472 480 512500 3946
rect 512656 3602 512684 6052
rect 513564 4072 513616 4078
rect 513564 4014 513616 4020
rect 512644 3596 512696 3602
rect 512644 3538 512696 3544
rect 513576 480 513604 4014
rect 513760 4010 513788 6052
rect 513748 4004 513800 4010
rect 513748 3946 513800 3952
rect 514864 3874 514892 6052
rect 515982 6038 516088 6066
rect 514852 3868 514904 3874
rect 514852 3810 514904 3816
rect 514760 3664 514812 3670
rect 514760 3606 514812 3612
rect 514772 480 514800 3606
rect 516060 3398 516088 6038
rect 515956 3392 516008 3398
rect 515956 3334 516008 3340
rect 516048 3392 516100 3398
rect 516048 3334 516100 3340
rect 515968 480 515996 3334
rect 517072 3194 517100 6052
rect 518176 3942 518204 6052
rect 517980 3936 518032 3942
rect 517980 3878 518032 3884
rect 518164 3936 518216 3942
rect 518164 3878 518216 3884
rect 517152 3324 517204 3330
rect 517152 3266 517204 3272
rect 517060 3188 517112 3194
rect 517060 3130 517112 3136
rect 517164 480 517192 3266
rect 468638 354 468750 480
rect 468312 326 468750 354
rect 468638 -960 468750 326
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 517992 354 518020 3878
rect 519280 3670 519308 6052
rect 520384 4078 520412 6052
rect 520372 4072 520424 4078
rect 520372 4014 520424 4020
rect 520740 3800 520792 3806
rect 520740 3742 520792 3748
rect 519268 3664 519320 3670
rect 519268 3606 519320 3612
rect 519544 3120 519596 3126
rect 519544 3062 519596 3068
rect 519556 480 519584 3062
rect 520752 480 520780 3742
rect 521488 3505 521516 6052
rect 521474 3496 521530 3505
rect 522592 3466 522620 6052
rect 523696 3534 523724 6052
rect 523040 3528 523092 3534
rect 523040 3470 523092 3476
rect 523684 3528 523736 3534
rect 523684 3470 523736 3476
rect 521474 3431 521530 3440
rect 521844 3460 521896 3466
rect 521844 3402 521896 3408
rect 522580 3460 522632 3466
rect 522580 3402 522632 3408
rect 521856 480 521884 3402
rect 523052 480 523080 3470
rect 524800 3330 524828 6052
rect 525904 4146 525932 6052
rect 525800 4140 525852 4146
rect 525800 4082 525852 4088
rect 525892 4140 525944 4146
rect 525892 4082 525944 4088
rect 524788 3324 524840 3330
rect 524788 3266 524840 3272
rect 525432 3256 525484 3262
rect 525432 3198 525484 3204
rect 524236 3052 524288 3058
rect 524236 2994 524288 3000
rect 524248 480 524276 2994
rect 525444 480 525472 3198
rect 525812 2854 525840 4082
rect 527008 3534 527036 6052
rect 528112 3738 528140 6052
rect 529216 3806 529244 6052
rect 530320 4010 530348 6052
rect 530124 4004 530176 4010
rect 530124 3946 530176 3952
rect 530308 4004 530360 4010
rect 530308 3946 530360 3952
rect 529204 3800 529256 3806
rect 529204 3742 529256 3748
rect 527824 3732 527876 3738
rect 527824 3674 527876 3680
rect 528100 3732 528152 3738
rect 528100 3674 528152 3680
rect 526720 3528 526772 3534
rect 526720 3470 526772 3476
rect 526996 3528 527048 3534
rect 526996 3470 527048 3476
rect 526732 3330 526760 3470
rect 526720 3324 526772 3330
rect 526720 3266 526772 3272
rect 525800 2848 525852 2854
rect 525800 2790 525852 2796
rect 526628 2848 526680 2854
rect 526628 2790 526680 2796
rect 526640 480 526668 2790
rect 527836 480 527864 3674
rect 529020 3596 529072 3602
rect 529020 3538 529072 3544
rect 529032 480 529060 3538
rect 530136 480 530164 3946
rect 531320 3868 531372 3874
rect 531320 3810 531372 3816
rect 531332 480 531360 3810
rect 531424 3126 531452 6052
rect 532542 6038 532648 6066
rect 532620 3398 532648 6038
rect 533632 3874 533660 6052
rect 534736 3942 534764 6052
rect 534540 3936 534592 3942
rect 534540 3878 534592 3884
rect 534724 3936 534776 3942
rect 534724 3878 534776 3884
rect 533620 3868 533672 3874
rect 533620 3810 533672 3816
rect 532516 3392 532568 3398
rect 532516 3334 532568 3340
rect 532608 3392 532660 3398
rect 532608 3334 532660 3340
rect 531412 3120 531464 3126
rect 531412 3062 531464 3068
rect 532528 480 532556 3334
rect 533712 3188 533764 3194
rect 533712 3130 533764 3136
rect 533724 480 533752 3130
rect 518318 354 518430 480
rect 517992 326 518430 354
rect 518318 -960 518430 326
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534552 354 534580 3878
rect 535840 3670 535868 6052
rect 536944 4078 536972 6052
rect 536840 4072 536892 4078
rect 536840 4014 536892 4020
rect 536932 4072 536984 4078
rect 536932 4014 536984 4020
rect 535828 3664 535880 3670
rect 535828 3606 535880 3612
rect 536104 3596 536156 3602
rect 536104 3538 536156 3544
rect 536116 480 536144 3538
rect 536852 2122 536880 4014
rect 538048 3369 538076 6052
rect 539152 3777 539180 6052
rect 539138 3768 539194 3777
rect 539138 3703 539194 3712
rect 538402 3496 538458 3505
rect 538402 3431 538458 3440
rect 539600 3460 539652 3466
rect 538034 3360 538090 3369
rect 538034 3295 538090 3304
rect 536852 2094 537248 2122
rect 537220 480 537248 2094
rect 538416 480 538444 3431
rect 539600 3402 539652 3408
rect 539612 480 539640 3402
rect 540256 3194 540284 6052
rect 540796 3324 540848 3330
rect 540796 3266 540848 3272
rect 540244 3188 540296 3194
rect 540244 3130 540296 3136
rect 540808 480 540836 3266
rect 541360 3058 541388 6052
rect 542464 3466 542492 6052
rect 543188 4140 543240 4146
rect 543188 4082 543240 4088
rect 542452 3460 542504 3466
rect 542452 3402 542504 3408
rect 541992 3256 542044 3262
rect 541992 3198 542044 3204
rect 541348 3052 541400 3058
rect 541348 2994 541400 3000
rect 542004 480 542032 3198
rect 543200 480 543228 4082
rect 543568 3602 543596 6052
rect 543556 3596 543608 3602
rect 543556 3538 543608 3544
rect 544672 3534 544700 6052
rect 545776 3738 545804 6052
rect 546684 3800 546736 3806
rect 546684 3742 546736 3748
rect 545488 3732 545540 3738
rect 545488 3674 545540 3680
rect 545764 3732 545816 3738
rect 545764 3674 545816 3680
rect 544384 3528 544436 3534
rect 544384 3470 544436 3476
rect 544660 3528 544712 3534
rect 544660 3470 544712 3476
rect 544396 480 544424 3470
rect 545500 480 545528 3674
rect 546696 480 546724 3742
rect 546880 3262 546908 6052
rect 547880 4004 547932 4010
rect 547880 3946 547932 3952
rect 546868 3256 546920 3262
rect 546868 3198 546920 3204
rect 547892 480 547920 3946
rect 547984 2990 548012 6052
rect 549088 4146 549116 6052
rect 549076 4140 549128 4146
rect 549076 4082 549128 4088
rect 550192 4010 550220 6052
rect 550180 4004 550232 4010
rect 550180 3946 550232 3952
rect 551296 3874 551324 6052
rect 551100 3868 551152 3874
rect 551100 3810 551152 3816
rect 551284 3868 551336 3874
rect 551284 3810 551336 3816
rect 550272 3392 550324 3398
rect 550272 3334 550324 3340
rect 549076 3120 549128 3126
rect 549076 3062 549128 3068
rect 547972 2984 548024 2990
rect 547972 2926 548024 2932
rect 549088 480 549116 3062
rect 550284 480 550312 3334
rect 534878 354 534990 480
rect 534552 326 534990 354
rect 534878 -960 534990 326
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551112 354 551140 3810
rect 552400 3641 552428 6052
rect 553504 3942 553532 6052
rect 552664 3936 552716 3942
rect 552664 3878 552716 3884
rect 553492 3936 553544 3942
rect 553492 3878 553544 3884
rect 552386 3632 552442 3641
rect 552386 3567 552442 3576
rect 552676 480 552704 3878
rect 553768 3664 553820 3670
rect 553768 3606 553820 3612
rect 553780 480 553808 3606
rect 554608 3398 554636 6052
rect 554964 4072 555016 4078
rect 554964 4014 555016 4020
rect 554596 3392 554648 3398
rect 554596 3334 554648 3340
rect 554976 480 555004 4014
rect 555712 3505 555740 6052
rect 556816 4078 556844 6052
rect 556804 4072 556856 4078
rect 556804 4014 556856 4020
rect 557920 3806 557948 6052
rect 557908 3800 557960 3806
rect 557354 3768 557410 3777
rect 557908 3742 557960 3748
rect 557354 3703 557410 3712
rect 555698 3496 555754 3505
rect 555698 3431 555754 3440
rect 556158 3360 556214 3369
rect 556158 3295 556214 3304
rect 556172 480 556200 3295
rect 557368 480 557396 3703
rect 559024 3670 559052 6052
rect 559012 3664 559064 3670
rect 559012 3606 559064 3612
rect 560128 3369 560156 6052
rect 561232 3466 561260 6052
rect 562336 3602 562364 6052
rect 562048 3596 562100 3602
rect 562048 3538 562100 3544
rect 562324 3596 562376 3602
rect 562324 3538 562376 3544
rect 560852 3460 560904 3466
rect 560852 3402 560904 3408
rect 561220 3460 561272 3466
rect 561220 3402 561272 3408
rect 560114 3360 560170 3369
rect 558552 3324 558604 3330
rect 560114 3295 560170 3304
rect 558552 3266 558604 3272
rect 558564 480 558592 3266
rect 559748 3188 559800 3194
rect 559748 3130 559800 3136
rect 559760 480 559788 3130
rect 560864 480 560892 3402
rect 562060 480 562088 3538
rect 563440 3534 563468 6052
rect 568028 4140 568080 4146
rect 568028 4082 568080 4088
rect 564440 3732 564492 3738
rect 564440 3674 564492 3680
rect 563244 3528 563296 3534
rect 563244 3470 563296 3476
rect 563428 3528 563480 3534
rect 563428 3470 563480 3476
rect 563256 480 563284 3470
rect 564452 480 564480 3674
rect 565636 3256 565688 3262
rect 565636 3198 565688 3204
rect 565648 480 565676 3198
rect 566832 3120 566884 3126
rect 566832 3062 566884 3068
rect 566844 480 566872 3062
rect 568040 480 568068 4082
rect 576308 4072 576360 4078
rect 576308 4014 576360 4020
rect 569132 4004 569184 4010
rect 569132 3946 569184 3952
rect 569144 480 569172 3946
rect 572720 3936 572772 3942
rect 572720 3878 572772 3884
rect 570328 3868 570380 3874
rect 570328 3810 570380 3816
rect 570340 480 570368 3810
rect 571522 3632 571578 3641
rect 571522 3567 571578 3576
rect 571536 480 571564 3567
rect 572732 480 572760 3878
rect 575110 3496 575166 3505
rect 575110 3431 575166 3440
rect 573916 3392 573968 3398
rect 573916 3334 573968 3340
rect 573928 480 573956 3334
rect 575124 480 575152 3431
rect 576320 480 576348 4014
rect 577412 3800 577464 3806
rect 577412 3742 577464 3748
rect 577424 480 577452 3742
rect 578608 3664 578660 3670
rect 578608 3606 578660 3612
rect 578620 480 578648 3606
rect 582196 3596 582248 3602
rect 582196 3538 582248 3544
rect 581000 3460 581052 3466
rect 581000 3402 581052 3408
rect 579802 3360 579858 3369
rect 579802 3295 579858 3304
rect 579816 480 579844 3295
rect 581012 480 581040 3402
rect 582208 480 582236 3538
rect 583392 3528 583444 3534
rect 583392 3470 583444 3476
rect 583404 480 583432 3470
rect 551438 354 551550 480
rect 551112 326 551550 354
rect 551438 -960 551550 326
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 697312 3478 697368
rect 578882 697176 578938 697232
rect 578882 685208 578938 685264
rect 3422 684392 3478 684448
rect 3606 684256 3662 684312
rect 580262 683848 580318 683904
rect 578330 672288 578386 672344
rect 3606 671744 3662 671800
rect 3422 671200 3478 671256
rect 580262 670656 580318 670712
rect 578514 659404 578516 659424
rect 578516 659404 578568 659424
rect 578568 659404 578570 659424
rect 578514 659368 578570 659404
rect 3422 659096 3478 659152
rect 3422 658144 3478 658200
rect 580262 657328 580318 657384
rect 3422 646448 3478 646504
rect 578330 646448 578386 646504
rect 3422 645088 3478 645144
rect 578882 644000 578938 644056
rect 3422 633800 3478 633856
rect 578882 633528 578938 633584
rect 3422 632032 3478 632088
rect 580262 630808 580318 630864
rect 3422 621152 3478 621208
rect 578330 620608 578386 620664
rect 3422 619112 3478 619168
rect 578882 617480 578938 617536
rect 3422 608504 3478 608560
rect 578882 607688 578938 607744
rect 3422 606056 3478 606112
rect 578882 604152 578938 604208
rect 3422 595856 3478 595912
rect 578882 594768 578938 594824
rect 3422 593000 3478 593056
rect 578882 590960 578938 591016
rect 3422 583208 3478 583264
rect 578882 581848 578938 581904
rect 3422 579944 3478 580000
rect 578882 577632 578938 577688
rect 3422 570560 3478 570616
rect 578882 568928 578938 568984
rect 3054 566888 3110 566944
rect 578882 564304 578938 564360
rect 3054 557912 3110 557968
rect 578882 556008 578938 556064
rect 3422 553832 3478 553888
rect 578882 551112 578938 551168
rect 3422 545264 3478 545320
rect 578882 543088 578938 543144
rect 2962 540776 3018 540832
rect 579526 537784 579582 537840
rect 2962 532616 3018 532672
rect 579526 530168 579582 530224
rect 2962 527856 3018 527912
rect 578882 524456 578938 524512
rect 2962 519968 3018 520024
rect 578882 517248 578938 517304
rect 3422 514800 3478 514856
rect 580538 511264 580594 511320
rect 3422 507320 3478 507376
rect 578238 504328 578294 504384
rect 3054 501744 3110 501800
rect 579526 497936 579582 497992
rect 3054 494672 3110 494728
rect 579526 491408 579582 491464
rect 2962 488688 3018 488744
rect 578882 484608 578938 484664
rect 2962 482024 3018 482080
rect 578882 478488 578938 478544
rect 3422 475632 3478 475688
rect 579802 471416 579858 471472
rect 3422 469376 3478 469432
rect 578238 465568 578294 465624
rect 2962 462576 3018 462632
rect 579526 458088 579582 458144
rect 2962 456728 3018 456784
rect 579526 452648 579582 452704
rect 3054 449520 3110 449576
rect 578882 444760 578938 444816
rect 3054 444080 3110 444136
rect 578882 439728 578938 439784
rect 3422 436600 3478 436656
rect 579526 431568 579582 431624
rect 3422 431432 3478 431488
rect 579526 426808 579582 426864
rect 2962 423544 3018 423600
rect 2962 418784 3018 418840
rect 579526 418240 579582 418296
rect 579526 413888 579582 413944
rect 3054 410488 3110 410544
rect 3054 406136 3110 406192
rect 580354 404912 580410 404968
rect 578238 400968 578294 401024
rect 2778 397432 2834 397488
rect 2778 393488 2834 393544
rect 579618 391720 579674 391776
rect 579526 388048 579582 388104
rect 3054 384376 3110 384432
rect 3054 380840 3110 380896
rect 579526 378392 579582 378448
rect 579526 375128 579582 375184
rect 3054 371320 3110 371376
rect 3054 368192 3110 368248
rect 580906 365064 580962 365120
rect 578330 362208 578386 362264
rect 3054 358400 3110 358456
rect 3054 355544 3110 355600
rect 579618 351872 579674 351928
rect 579526 349288 579582 349344
rect 3054 345344 3110 345400
rect 3054 342896 3110 342952
rect 579618 338544 579674 338600
rect 579526 336368 579582 336424
rect 3054 332288 3110 332344
rect 3054 330248 3110 330304
rect 579618 325216 579674 325272
rect 579526 323448 579582 323504
rect 3054 319232 3110 319288
rect 3054 317600 3110 317656
rect 579618 312024 579674 312080
rect 579526 310528 579582 310584
rect 3054 306176 3110 306232
rect 3054 304952 3110 305008
rect 579618 298696 579674 298752
rect 579526 297608 579582 297664
rect 3054 293120 3110 293176
rect 3054 292304 3110 292360
rect 3054 229064 3110 229120
rect 3054 227976 3110 228032
rect 578514 220088 578570 220144
rect 580906 219000 580962 219056
rect 3054 216416 3110 216472
rect 3054 214920 3110 214976
rect 579526 207168 579582 207224
rect 579618 205672 579674 205728
rect 3054 203768 3110 203824
rect 3054 201864 3110 201920
rect 579526 194248 579582 194304
rect 579618 192480 579674 192536
rect 2962 191120 3018 191176
rect 2962 188808 3018 188864
rect 578330 181348 578386 181384
rect 578330 181328 578332 181348
rect 578332 181328 578384 181348
rect 578384 181328 578386 181348
rect 580538 179152 580594 179208
rect 2962 178472 3018 178528
rect 2962 175888 3018 175944
rect 579526 168408 579582 168464
rect 3054 165824 3110 165880
rect 579618 165824 579674 165880
rect 3054 162832 3110 162888
rect 579526 155488 579582 155544
rect 3054 153176 3110 153232
rect 579618 152632 579674 152688
rect 3054 149776 3110 149832
rect 578790 142588 578846 142624
rect 578790 142568 578792 142588
rect 578792 142568 578844 142588
rect 578844 142568 578846 142588
rect 3054 140528 3110 140584
rect 580722 139304 580778 139360
rect 3054 136720 3110 136776
rect 579526 129648 579582 129704
rect 3054 127880 3110 127936
rect 579618 125976 579674 126032
rect 3054 123664 3110 123720
rect 578330 116748 578386 116784
rect 578330 116728 578332 116748
rect 578332 116728 578384 116748
rect 578384 116728 578386 116748
rect 2962 115232 3018 115288
rect 580262 112784 580318 112840
rect 2962 110608 3018 110664
rect 579526 103808 579582 103864
rect 3054 102584 3110 102640
rect 579802 99456 579858 99512
rect 3054 97552 3110 97608
rect 579526 90888 579582 90944
rect 3054 89936 3110 89992
rect 579618 86128 579674 86184
rect 3054 84632 3110 84688
rect 578882 77968 578938 78024
rect 3422 77288 3478 77344
rect 578882 72936 578938 72992
rect 3422 71576 3478 71632
rect 578238 65048 578294 65104
rect 3054 64640 3110 64696
rect 580814 59608 580870 59664
rect 3054 58520 3110 58576
rect 579526 52128 579582 52184
rect 3422 51992 3478 52048
rect 579526 46280 579582 46336
rect 3422 45464 3478 45520
rect 3422 39344 3478 39400
rect 578882 39208 578938 39264
rect 578882 33088 578938 33144
rect 3422 32408 3478 32464
rect 2962 26696 3018 26752
rect 578238 26288 578294 26344
rect 580630 19760 580686 19816
rect 2962 19352 3018 19408
rect 3422 14048 3478 14104
rect 578882 13368 578938 13424
rect 578882 6568 578938 6624
rect 3422 6432 3478 6488
rect 5262 3304 5318 3360
rect 20626 3440 20682 3496
rect 23570 3304 23626 3360
rect 28906 3304 28962 3360
rect 37922 3440 37978 3496
rect 45650 3304 45706 3360
rect 521474 3440 521530 3496
rect 539138 3712 539194 3768
rect 538402 3440 538458 3496
rect 538034 3304 538090 3360
rect 552386 3576 552442 3632
rect 557354 3712 557410 3768
rect 555698 3440 555754 3496
rect 556158 3304 556214 3360
rect 560114 3304 560170 3360
rect 571522 3576 571578 3632
rect 575110 3440 575166 3496
rect 579802 3304 579858 3360
<< metal3 >>
rect -960 697370 480 697460
rect 3417 697370 3483 697373
rect -960 697368 3483 697370
rect -960 697312 3422 697368
rect 3478 697312 3483 697368
rect -960 697310 3483 697312
rect -960 697220 480 697310
rect 3417 697307 3483 697310
rect 578877 697234 578943 697237
rect 583520 697234 584960 697324
rect 578877 697232 584960 697234
rect 578877 697176 578882 697232
rect 578938 697176 584960 697232
rect 578877 697174 584960 697176
rect 578877 697171 578943 697174
rect 583520 697084 584960 697174
rect 578877 685266 578943 685269
rect 576748 685264 578943 685266
rect 576748 685208 578882 685264
rect 578938 685208 578943 685264
rect 576748 685206 578943 685208
rect 578877 685203 578943 685206
rect 3417 684450 3483 684453
rect 3417 684448 6164 684450
rect -960 684314 480 684404
rect 3417 684392 3422 684448
rect 3478 684392 6164 684448
rect 3417 684390 6164 684392
rect 3417 684387 3483 684390
rect 3601 684314 3667 684317
rect -960 684312 3667 684314
rect -960 684256 3606 684312
rect 3662 684256 3667 684312
rect -960 684254 3667 684256
rect -960 684164 480 684254
rect 3601 684251 3667 684254
rect 580257 683906 580323 683909
rect 583520 683906 584960 683996
rect 580257 683904 584960 683906
rect 580257 683848 580262 683904
rect 580318 683848 584960 683904
rect 580257 683846 584960 683848
rect 580257 683843 580323 683846
rect 583520 683756 584960 683846
rect 578325 672346 578391 672349
rect 576748 672344 578391 672346
rect 576748 672288 578330 672344
rect 578386 672288 578391 672344
rect 576748 672286 578391 672288
rect 578325 672283 578391 672286
rect 3601 671802 3667 671805
rect 3601 671800 6164 671802
rect 3601 671744 3606 671800
rect 3662 671744 6164 671800
rect 3601 671742 6164 671744
rect 3601 671739 3667 671742
rect -960 671258 480 671348
rect 3417 671258 3483 671261
rect -960 671256 3483 671258
rect -960 671200 3422 671256
rect 3478 671200 3483 671256
rect -960 671198 3483 671200
rect -960 671108 480 671198
rect 3417 671195 3483 671198
rect 580257 670714 580323 670717
rect 583520 670714 584960 670804
rect 580257 670712 584960 670714
rect 580257 670656 580262 670712
rect 580318 670656 584960 670712
rect 580257 670654 584960 670656
rect 580257 670651 580323 670654
rect 583520 670564 584960 670654
rect 578509 659426 578575 659429
rect 576748 659424 578575 659426
rect 576748 659368 578514 659424
rect 578570 659368 578575 659424
rect 576748 659366 578575 659368
rect 578509 659363 578575 659366
rect 3417 659154 3483 659157
rect 3417 659152 6164 659154
rect 3417 659096 3422 659152
rect 3478 659096 6164 659152
rect 3417 659094 6164 659096
rect 3417 659091 3483 659094
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 580257 657386 580323 657389
rect 583520 657386 584960 657476
rect 580257 657384 584960 657386
rect 580257 657328 580262 657384
rect 580318 657328 584960 657384
rect 580257 657326 584960 657328
rect 580257 657323 580323 657326
rect 583520 657236 584960 657326
rect 3417 646506 3483 646509
rect 578325 646506 578391 646509
rect 3417 646504 6164 646506
rect 3417 646448 3422 646504
rect 3478 646448 6164 646504
rect 3417 646446 6164 646448
rect 576748 646504 578391 646506
rect 576748 646448 578330 646504
rect 578386 646448 578391 646504
rect 576748 646446 578391 646448
rect 3417 646443 3483 646446
rect 578325 646443 578391 646446
rect -960 645146 480 645236
rect 3417 645146 3483 645149
rect -960 645144 3483 645146
rect -960 645088 3422 645144
rect 3478 645088 3483 645144
rect -960 645086 3483 645088
rect -960 644996 480 645086
rect 3417 645083 3483 645086
rect 578877 644058 578943 644061
rect 583520 644058 584960 644148
rect 578877 644056 584960 644058
rect 578877 644000 578882 644056
rect 578938 644000 584960 644056
rect 578877 643998 584960 644000
rect 578877 643995 578943 643998
rect 583520 643908 584960 643998
rect 3417 633858 3483 633861
rect 3417 633856 6164 633858
rect 3417 633800 3422 633856
rect 3478 633800 6164 633856
rect 3417 633798 6164 633800
rect 3417 633795 3483 633798
rect 578877 633586 578943 633589
rect 576748 633584 578943 633586
rect 576748 633528 578882 633584
rect 578938 633528 578943 633584
rect 576748 633526 578943 633528
rect 578877 633523 578943 633526
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 580257 630866 580323 630869
rect 583520 630866 584960 630956
rect 580257 630864 584960 630866
rect 580257 630808 580262 630864
rect 580318 630808 584960 630864
rect 580257 630806 584960 630808
rect 580257 630803 580323 630806
rect 583520 630716 584960 630806
rect 3417 621210 3483 621213
rect 3417 621208 6164 621210
rect 3417 621152 3422 621208
rect 3478 621152 6164 621208
rect 3417 621150 6164 621152
rect 3417 621147 3483 621150
rect 578325 620666 578391 620669
rect 576748 620664 578391 620666
rect 576748 620608 578330 620664
rect 578386 620608 578391 620664
rect 576748 620606 578391 620608
rect 578325 620603 578391 620606
rect -960 619170 480 619260
rect 3417 619170 3483 619173
rect -960 619168 3483 619170
rect -960 619112 3422 619168
rect 3478 619112 3483 619168
rect -960 619110 3483 619112
rect -960 619020 480 619110
rect 3417 619107 3483 619110
rect 578877 617538 578943 617541
rect 583520 617538 584960 617628
rect 578877 617536 584960 617538
rect 578877 617480 578882 617536
rect 578938 617480 584960 617536
rect 578877 617478 584960 617480
rect 578877 617475 578943 617478
rect 583520 617388 584960 617478
rect 3417 608562 3483 608565
rect 3417 608560 6164 608562
rect 3417 608504 3422 608560
rect 3478 608504 6164 608560
rect 3417 608502 6164 608504
rect 3417 608499 3483 608502
rect 578877 607746 578943 607749
rect 576748 607744 578943 607746
rect 576748 607688 578882 607744
rect 578938 607688 578943 607744
rect 576748 607686 578943 607688
rect 578877 607683 578943 607686
rect -960 606114 480 606204
rect 3417 606114 3483 606117
rect -960 606112 3483 606114
rect -960 606056 3422 606112
rect 3478 606056 3483 606112
rect -960 606054 3483 606056
rect -960 605964 480 606054
rect 3417 606051 3483 606054
rect 578877 604210 578943 604213
rect 583520 604210 584960 604300
rect 578877 604208 584960 604210
rect 578877 604152 578882 604208
rect 578938 604152 584960 604208
rect 578877 604150 584960 604152
rect 578877 604147 578943 604150
rect 583520 604060 584960 604150
rect 3417 595914 3483 595917
rect 3417 595912 6164 595914
rect 3417 595856 3422 595912
rect 3478 595856 6164 595912
rect 3417 595854 6164 595856
rect 3417 595851 3483 595854
rect 578877 594826 578943 594829
rect 576748 594824 578943 594826
rect 576748 594768 578882 594824
rect 578938 594768 578943 594824
rect 576748 594766 578943 594768
rect 578877 594763 578943 594766
rect -960 593058 480 593148
rect 3417 593058 3483 593061
rect -960 593056 3483 593058
rect -960 593000 3422 593056
rect 3478 593000 3483 593056
rect -960 592998 3483 593000
rect -960 592908 480 592998
rect 3417 592995 3483 592998
rect 578877 591018 578943 591021
rect 583520 591018 584960 591108
rect 578877 591016 584960 591018
rect 578877 590960 578882 591016
rect 578938 590960 584960 591016
rect 578877 590958 584960 590960
rect 578877 590955 578943 590958
rect 583520 590868 584960 590958
rect 3417 583266 3483 583269
rect 3417 583264 6164 583266
rect 3417 583208 3422 583264
rect 3478 583208 6164 583264
rect 3417 583206 6164 583208
rect 3417 583203 3483 583206
rect 578877 581906 578943 581909
rect 576748 581904 578943 581906
rect 576748 581848 578882 581904
rect 578938 581848 578943 581904
rect 576748 581846 578943 581848
rect 578877 581843 578943 581846
rect -960 580002 480 580092
rect 3417 580002 3483 580005
rect -960 580000 3483 580002
rect -960 579944 3422 580000
rect 3478 579944 3483 580000
rect -960 579942 3483 579944
rect -960 579852 480 579942
rect 3417 579939 3483 579942
rect 578877 577690 578943 577693
rect 583520 577690 584960 577780
rect 578877 577688 584960 577690
rect 578877 577632 578882 577688
rect 578938 577632 584960 577688
rect 578877 577630 584960 577632
rect 578877 577627 578943 577630
rect 583520 577540 584960 577630
rect 3417 570618 3483 570621
rect 3417 570616 6164 570618
rect 3417 570560 3422 570616
rect 3478 570560 6164 570616
rect 3417 570558 6164 570560
rect 3417 570555 3483 570558
rect 578877 568986 578943 568989
rect 576748 568984 578943 568986
rect 576748 568928 578882 568984
rect 578938 568928 578943 568984
rect 576748 568926 578943 568928
rect 578877 568923 578943 568926
rect -960 566946 480 567036
rect 3049 566946 3115 566949
rect -960 566944 3115 566946
rect -960 566888 3054 566944
rect 3110 566888 3115 566944
rect -960 566886 3115 566888
rect -960 566796 480 566886
rect 3049 566883 3115 566886
rect 578877 564362 578943 564365
rect 583520 564362 584960 564452
rect 578877 564360 584960 564362
rect 578877 564304 578882 564360
rect 578938 564304 584960 564360
rect 578877 564302 584960 564304
rect 578877 564299 578943 564302
rect 583520 564212 584960 564302
rect 3049 557970 3115 557973
rect 3049 557968 6164 557970
rect 3049 557912 3054 557968
rect 3110 557912 6164 557968
rect 3049 557910 6164 557912
rect 3049 557907 3115 557910
rect 578877 556066 578943 556069
rect 576748 556064 578943 556066
rect 576748 556008 578882 556064
rect 578938 556008 578943 556064
rect 576748 556006 578943 556008
rect 578877 556003 578943 556006
rect -960 553890 480 553980
rect 3417 553890 3483 553893
rect -960 553888 3483 553890
rect -960 553832 3422 553888
rect 3478 553832 3483 553888
rect -960 553830 3483 553832
rect -960 553740 480 553830
rect 3417 553827 3483 553830
rect 578877 551170 578943 551173
rect 583520 551170 584960 551260
rect 578877 551168 584960 551170
rect 578877 551112 578882 551168
rect 578938 551112 584960 551168
rect 578877 551110 584960 551112
rect 578877 551107 578943 551110
rect 583520 551020 584960 551110
rect 3417 545322 3483 545325
rect 3417 545320 6164 545322
rect 3417 545264 3422 545320
rect 3478 545264 6164 545320
rect 3417 545262 6164 545264
rect 3417 545259 3483 545262
rect 578877 543146 578943 543149
rect 576748 543144 578943 543146
rect 576748 543088 578882 543144
rect 578938 543088 578943 543144
rect 576748 543086 578943 543088
rect 578877 543083 578943 543086
rect -960 540834 480 540924
rect 2957 540834 3023 540837
rect -960 540832 3023 540834
rect -960 540776 2962 540832
rect 3018 540776 3023 540832
rect -960 540774 3023 540776
rect -960 540684 480 540774
rect 2957 540771 3023 540774
rect 579521 537842 579587 537845
rect 583520 537842 584960 537932
rect 579521 537840 584960 537842
rect 579521 537784 579526 537840
rect 579582 537784 584960 537840
rect 579521 537782 584960 537784
rect 579521 537779 579587 537782
rect 583520 537692 584960 537782
rect 2957 532674 3023 532677
rect 2957 532672 6164 532674
rect 2957 532616 2962 532672
rect 3018 532616 6164 532672
rect 2957 532614 6164 532616
rect 2957 532611 3023 532614
rect 579521 530226 579587 530229
rect 576748 530224 579587 530226
rect 576748 530168 579526 530224
rect 579582 530168 579587 530224
rect 576748 530166 579587 530168
rect 579521 530163 579587 530166
rect -960 527914 480 528004
rect 2957 527914 3023 527917
rect -960 527912 3023 527914
rect -960 527856 2962 527912
rect 3018 527856 3023 527912
rect -960 527854 3023 527856
rect -960 527764 480 527854
rect 2957 527851 3023 527854
rect 578877 524514 578943 524517
rect 583520 524514 584960 524604
rect 578877 524512 584960 524514
rect 578877 524456 578882 524512
rect 578938 524456 584960 524512
rect 578877 524454 584960 524456
rect 578877 524451 578943 524454
rect 583520 524364 584960 524454
rect 2957 520026 3023 520029
rect 2957 520024 6164 520026
rect 2957 519968 2962 520024
rect 3018 519968 6164 520024
rect 2957 519966 6164 519968
rect 2957 519963 3023 519966
rect 578877 517306 578943 517309
rect 576748 517304 578943 517306
rect 576748 517248 578882 517304
rect 578938 517248 578943 517304
rect 576748 517246 578943 517248
rect 578877 517243 578943 517246
rect -960 514858 480 514948
rect 3417 514858 3483 514861
rect -960 514856 3483 514858
rect -960 514800 3422 514856
rect 3478 514800 3483 514856
rect -960 514798 3483 514800
rect -960 514708 480 514798
rect 3417 514795 3483 514798
rect 580533 511322 580599 511325
rect 583520 511322 584960 511412
rect 580533 511320 584960 511322
rect 580533 511264 580538 511320
rect 580594 511264 584960 511320
rect 580533 511262 584960 511264
rect 580533 511259 580599 511262
rect 583520 511172 584960 511262
rect 3417 507378 3483 507381
rect 3417 507376 6164 507378
rect 3417 507320 3422 507376
rect 3478 507320 6164 507376
rect 3417 507318 6164 507320
rect 3417 507315 3483 507318
rect 578233 504386 578299 504389
rect 576748 504384 578299 504386
rect 576748 504328 578238 504384
rect 578294 504328 578299 504384
rect 576748 504326 578299 504328
rect 578233 504323 578299 504326
rect -960 501802 480 501892
rect 3049 501802 3115 501805
rect -960 501800 3115 501802
rect -960 501744 3054 501800
rect 3110 501744 3115 501800
rect -960 501742 3115 501744
rect -960 501652 480 501742
rect 3049 501739 3115 501742
rect 579521 497994 579587 497997
rect 583520 497994 584960 498084
rect 579521 497992 584960 497994
rect 579521 497936 579526 497992
rect 579582 497936 584960 497992
rect 579521 497934 584960 497936
rect 579521 497931 579587 497934
rect 583520 497844 584960 497934
rect 3049 494730 3115 494733
rect 3049 494728 6164 494730
rect 3049 494672 3054 494728
rect 3110 494672 6164 494728
rect 3049 494670 6164 494672
rect 3049 494667 3115 494670
rect 579521 491466 579587 491469
rect 576748 491464 579587 491466
rect 576748 491408 579526 491464
rect 579582 491408 579587 491464
rect 576748 491406 579587 491408
rect 579521 491403 579587 491406
rect -960 488746 480 488836
rect 2957 488746 3023 488749
rect -960 488744 3023 488746
rect -960 488688 2962 488744
rect 3018 488688 3023 488744
rect -960 488686 3023 488688
rect -960 488596 480 488686
rect 2957 488683 3023 488686
rect 578877 484666 578943 484669
rect 583520 484666 584960 484756
rect 578877 484664 584960 484666
rect 578877 484608 578882 484664
rect 578938 484608 584960 484664
rect 578877 484606 584960 484608
rect 578877 484603 578943 484606
rect 583520 484516 584960 484606
rect 2957 482082 3023 482085
rect 2957 482080 6164 482082
rect 2957 482024 2962 482080
rect 3018 482024 6164 482080
rect 2957 482022 6164 482024
rect 2957 482019 3023 482022
rect 578877 478546 578943 478549
rect 576748 478544 578943 478546
rect 576748 478488 578882 478544
rect 578938 478488 578943 478544
rect 576748 478486 578943 478488
rect 578877 478483 578943 478486
rect -960 475690 480 475780
rect 3417 475690 3483 475693
rect -960 475688 3483 475690
rect -960 475632 3422 475688
rect 3478 475632 3483 475688
rect -960 475630 3483 475632
rect -960 475540 480 475630
rect 3417 475627 3483 475630
rect 579797 471474 579863 471477
rect 583520 471474 584960 471564
rect 579797 471472 584960 471474
rect 579797 471416 579802 471472
rect 579858 471416 584960 471472
rect 579797 471414 584960 471416
rect 579797 471411 579863 471414
rect 583520 471324 584960 471414
rect 3417 469434 3483 469437
rect 3417 469432 6164 469434
rect 3417 469376 3422 469432
rect 3478 469376 6164 469432
rect 3417 469374 6164 469376
rect 3417 469371 3483 469374
rect 578233 465626 578299 465629
rect 576748 465624 578299 465626
rect 576748 465568 578238 465624
rect 578294 465568 578299 465624
rect 576748 465566 578299 465568
rect 578233 465563 578299 465566
rect -960 462634 480 462724
rect 2957 462634 3023 462637
rect -960 462632 3023 462634
rect -960 462576 2962 462632
rect 3018 462576 3023 462632
rect -960 462574 3023 462576
rect -960 462484 480 462574
rect 2957 462571 3023 462574
rect 579521 458146 579587 458149
rect 583520 458146 584960 458236
rect 579521 458144 584960 458146
rect 579521 458088 579526 458144
rect 579582 458088 584960 458144
rect 579521 458086 584960 458088
rect 579521 458083 579587 458086
rect 583520 457996 584960 458086
rect 2957 456786 3023 456789
rect 2957 456784 6164 456786
rect 2957 456728 2962 456784
rect 3018 456728 6164 456784
rect 2957 456726 6164 456728
rect 2957 456723 3023 456726
rect 579521 452706 579587 452709
rect 576748 452704 579587 452706
rect 576748 452648 579526 452704
rect 579582 452648 579587 452704
rect 576748 452646 579587 452648
rect 579521 452643 579587 452646
rect -960 449578 480 449668
rect 3049 449578 3115 449581
rect -960 449576 3115 449578
rect -960 449520 3054 449576
rect 3110 449520 3115 449576
rect -960 449518 3115 449520
rect -960 449428 480 449518
rect 3049 449515 3115 449518
rect 578877 444818 578943 444821
rect 583520 444818 584960 444908
rect 578877 444816 584960 444818
rect 578877 444760 578882 444816
rect 578938 444760 584960 444816
rect 578877 444758 584960 444760
rect 578877 444755 578943 444758
rect 583520 444668 584960 444758
rect 3049 444138 3115 444141
rect 3049 444136 6164 444138
rect 3049 444080 3054 444136
rect 3110 444080 6164 444136
rect 3049 444078 6164 444080
rect 3049 444075 3115 444078
rect 578877 439786 578943 439789
rect 576748 439784 578943 439786
rect 576748 439728 578882 439784
rect 578938 439728 578943 439784
rect 576748 439726 578943 439728
rect 578877 439723 578943 439726
rect -960 436658 480 436748
rect 3417 436658 3483 436661
rect -960 436656 3483 436658
rect -960 436600 3422 436656
rect 3478 436600 3483 436656
rect -960 436598 3483 436600
rect -960 436508 480 436598
rect 3417 436595 3483 436598
rect 579521 431626 579587 431629
rect 583520 431626 584960 431716
rect 579521 431624 584960 431626
rect 579521 431568 579526 431624
rect 579582 431568 584960 431624
rect 579521 431566 584960 431568
rect 579521 431563 579587 431566
rect 3417 431490 3483 431493
rect 3417 431488 6164 431490
rect 3417 431432 3422 431488
rect 3478 431432 6164 431488
rect 583520 431476 584960 431566
rect 3417 431430 6164 431432
rect 3417 431427 3483 431430
rect 579521 426866 579587 426869
rect 576748 426864 579587 426866
rect 576748 426808 579526 426864
rect 579582 426808 579587 426864
rect 576748 426806 579587 426808
rect 579521 426803 579587 426806
rect -960 423602 480 423692
rect 2957 423602 3023 423605
rect -960 423600 3023 423602
rect -960 423544 2962 423600
rect 3018 423544 3023 423600
rect -960 423542 3023 423544
rect -960 423452 480 423542
rect 2957 423539 3023 423542
rect 2957 418842 3023 418845
rect 2957 418840 6164 418842
rect 2957 418784 2962 418840
rect 3018 418784 6164 418840
rect 2957 418782 6164 418784
rect 2957 418779 3023 418782
rect 579521 418298 579587 418301
rect 583520 418298 584960 418388
rect 579521 418296 584960 418298
rect 579521 418240 579526 418296
rect 579582 418240 584960 418296
rect 579521 418238 584960 418240
rect 579521 418235 579587 418238
rect 583520 418148 584960 418238
rect 579521 413946 579587 413949
rect 576748 413944 579587 413946
rect 576748 413888 579526 413944
rect 579582 413888 579587 413944
rect 576748 413886 579587 413888
rect 579521 413883 579587 413886
rect -960 410546 480 410636
rect 3049 410546 3115 410549
rect -960 410544 3115 410546
rect -960 410488 3054 410544
rect 3110 410488 3115 410544
rect -960 410486 3115 410488
rect -960 410396 480 410486
rect 3049 410483 3115 410486
rect 3049 406194 3115 406197
rect 3049 406192 6164 406194
rect 3049 406136 3054 406192
rect 3110 406136 6164 406192
rect 3049 406134 6164 406136
rect 3049 406131 3115 406134
rect 580349 404970 580415 404973
rect 583520 404970 584960 405060
rect 580349 404968 584960 404970
rect 580349 404912 580354 404968
rect 580410 404912 584960 404968
rect 580349 404910 584960 404912
rect 580349 404907 580415 404910
rect 583520 404820 584960 404910
rect 578233 401026 578299 401029
rect 576748 401024 578299 401026
rect 576748 400968 578238 401024
rect 578294 400968 578299 401024
rect 576748 400966 578299 400968
rect 578233 400963 578299 400966
rect -960 397490 480 397580
rect 2773 397490 2839 397493
rect -960 397488 2839 397490
rect -960 397432 2778 397488
rect 2834 397432 2839 397488
rect -960 397430 2839 397432
rect -960 397340 480 397430
rect 2773 397427 2839 397430
rect 2773 393546 2839 393549
rect 2773 393544 6164 393546
rect 2773 393488 2778 393544
rect 2834 393488 6164 393544
rect 2773 393486 6164 393488
rect 2773 393483 2839 393486
rect 579613 391778 579679 391781
rect 583520 391778 584960 391868
rect 579613 391776 584960 391778
rect 579613 391720 579618 391776
rect 579674 391720 584960 391776
rect 579613 391718 584960 391720
rect 579613 391715 579679 391718
rect 583520 391628 584960 391718
rect 579521 388106 579587 388109
rect 576748 388104 579587 388106
rect 576748 388048 579526 388104
rect 579582 388048 579587 388104
rect 576748 388046 579587 388048
rect 579521 388043 579587 388046
rect -960 384434 480 384524
rect 3049 384434 3115 384437
rect -960 384432 3115 384434
rect -960 384376 3054 384432
rect 3110 384376 3115 384432
rect -960 384374 3115 384376
rect -960 384284 480 384374
rect 3049 384371 3115 384374
rect 3049 380898 3115 380901
rect 3049 380896 6164 380898
rect 3049 380840 3054 380896
rect 3110 380840 6164 380896
rect 3049 380838 6164 380840
rect 3049 380835 3115 380838
rect 579521 378450 579587 378453
rect 583520 378450 584960 378540
rect 579521 378448 584960 378450
rect 579521 378392 579526 378448
rect 579582 378392 584960 378448
rect 579521 378390 584960 378392
rect 579521 378387 579587 378390
rect 583520 378300 584960 378390
rect 579521 375186 579587 375189
rect 576748 375184 579587 375186
rect 576748 375128 579526 375184
rect 579582 375128 579587 375184
rect 576748 375126 579587 375128
rect 579521 375123 579587 375126
rect -960 371378 480 371468
rect 3049 371378 3115 371381
rect -960 371376 3115 371378
rect -960 371320 3054 371376
rect 3110 371320 3115 371376
rect -960 371318 3115 371320
rect -960 371228 480 371318
rect 3049 371315 3115 371318
rect 3049 368250 3115 368253
rect 3049 368248 6164 368250
rect 3049 368192 3054 368248
rect 3110 368192 6164 368248
rect 3049 368190 6164 368192
rect 3049 368187 3115 368190
rect 580901 365122 580967 365125
rect 583520 365122 584960 365212
rect 580901 365120 584960 365122
rect 580901 365064 580906 365120
rect 580962 365064 584960 365120
rect 580901 365062 584960 365064
rect 580901 365059 580967 365062
rect 583520 364972 584960 365062
rect 578325 362266 578391 362269
rect 576748 362264 578391 362266
rect 576748 362208 578330 362264
rect 578386 362208 578391 362264
rect 576748 362206 578391 362208
rect 578325 362203 578391 362206
rect -960 358458 480 358548
rect 3049 358458 3115 358461
rect -960 358456 3115 358458
rect -960 358400 3054 358456
rect 3110 358400 3115 358456
rect -960 358398 3115 358400
rect -960 358308 480 358398
rect 3049 358395 3115 358398
rect 3049 355602 3115 355605
rect 3049 355600 6164 355602
rect 3049 355544 3054 355600
rect 3110 355544 6164 355600
rect 3049 355542 6164 355544
rect 3049 355539 3115 355542
rect 579613 351930 579679 351933
rect 583520 351930 584960 352020
rect 579613 351928 584960 351930
rect 579613 351872 579618 351928
rect 579674 351872 584960 351928
rect 579613 351870 584960 351872
rect 579613 351867 579679 351870
rect 583520 351780 584960 351870
rect 579521 349346 579587 349349
rect 576748 349344 579587 349346
rect 576748 349288 579526 349344
rect 579582 349288 579587 349344
rect 576748 349286 579587 349288
rect 579521 349283 579587 349286
rect -960 345402 480 345492
rect 3049 345402 3115 345405
rect -960 345400 3115 345402
rect -960 345344 3054 345400
rect 3110 345344 3115 345400
rect -960 345342 3115 345344
rect -960 345252 480 345342
rect 3049 345339 3115 345342
rect 3049 342954 3115 342957
rect 3049 342952 6164 342954
rect 3049 342896 3054 342952
rect 3110 342896 6164 342952
rect 3049 342894 6164 342896
rect 3049 342891 3115 342894
rect 579613 338602 579679 338605
rect 583520 338602 584960 338692
rect 579613 338600 584960 338602
rect 579613 338544 579618 338600
rect 579674 338544 584960 338600
rect 579613 338542 584960 338544
rect 579613 338539 579679 338542
rect 583520 338452 584960 338542
rect 579521 336426 579587 336429
rect 576748 336424 579587 336426
rect 576748 336368 579526 336424
rect 579582 336368 579587 336424
rect 576748 336366 579587 336368
rect 579521 336363 579587 336366
rect -960 332346 480 332436
rect 3049 332346 3115 332349
rect -960 332344 3115 332346
rect -960 332288 3054 332344
rect 3110 332288 3115 332344
rect -960 332286 3115 332288
rect -960 332196 480 332286
rect 3049 332283 3115 332286
rect 3049 330306 3115 330309
rect 3049 330304 6164 330306
rect 3049 330248 3054 330304
rect 3110 330248 6164 330304
rect 3049 330246 6164 330248
rect 3049 330243 3115 330246
rect 579613 325274 579679 325277
rect 583520 325274 584960 325364
rect 579613 325272 584960 325274
rect 579613 325216 579618 325272
rect 579674 325216 584960 325272
rect 579613 325214 584960 325216
rect 579613 325211 579679 325214
rect 583520 325124 584960 325214
rect 579521 323506 579587 323509
rect 576748 323504 579587 323506
rect 576748 323448 579526 323504
rect 579582 323448 579587 323504
rect 576748 323446 579587 323448
rect 579521 323443 579587 323446
rect -960 319290 480 319380
rect 3049 319290 3115 319293
rect -960 319288 3115 319290
rect -960 319232 3054 319288
rect 3110 319232 3115 319288
rect -960 319230 3115 319232
rect -960 319140 480 319230
rect 3049 319227 3115 319230
rect 3049 317658 3115 317661
rect 3049 317656 6164 317658
rect 3049 317600 3054 317656
rect 3110 317600 6164 317656
rect 3049 317598 6164 317600
rect 3049 317595 3115 317598
rect 579613 312082 579679 312085
rect 583520 312082 584960 312172
rect 579613 312080 584960 312082
rect 579613 312024 579618 312080
rect 579674 312024 584960 312080
rect 579613 312022 584960 312024
rect 579613 312019 579679 312022
rect 583520 311932 584960 312022
rect 579521 310586 579587 310589
rect 576748 310584 579587 310586
rect 576748 310528 579526 310584
rect 579582 310528 579587 310584
rect 576748 310526 579587 310528
rect 579521 310523 579587 310526
rect -960 306234 480 306324
rect 3049 306234 3115 306237
rect -960 306232 3115 306234
rect -960 306176 3054 306232
rect 3110 306176 3115 306232
rect -960 306174 3115 306176
rect -960 306084 480 306174
rect 3049 306171 3115 306174
rect 3049 305010 3115 305013
rect 3049 305008 6164 305010
rect 3049 304952 3054 305008
rect 3110 304952 6164 305008
rect 3049 304950 6164 304952
rect 3049 304947 3115 304950
rect 579613 298754 579679 298757
rect 583520 298754 584960 298844
rect 579613 298752 584960 298754
rect 579613 298696 579618 298752
rect 579674 298696 584960 298752
rect 579613 298694 584960 298696
rect 579613 298691 579679 298694
rect 583520 298604 584960 298694
rect 579521 297666 579587 297669
rect 576748 297664 579587 297666
rect 576748 297608 579526 297664
rect 579582 297608 579587 297664
rect 576748 297606 579587 297608
rect 579521 297603 579587 297606
rect -960 293178 480 293268
rect 3049 293178 3115 293181
rect -960 293176 3115 293178
rect -960 293120 3054 293176
rect 3110 293120 3115 293176
rect -960 293118 3115 293120
rect -960 293028 480 293118
rect 3049 293115 3115 293118
rect 3049 292362 3115 292365
rect 3049 292360 6164 292362
rect 3049 292304 3054 292360
rect 3110 292304 6164 292360
rect 3049 292302 6164 292304
rect 3049 292299 3115 292302
rect 583520 285426 584960 285516
rect 583342 285366 584960 285426
rect 583342 285290 583402 285366
rect 583520 285290 584960 285366
rect 583342 285276 584960 285290
rect 583342 285230 583586 285276
rect 583526 284746 583586 285230
rect 576748 284686 583586 284746
rect -960 280122 480 280212
rect -960 280062 6194 280122
rect -960 279972 480 280062
rect 6134 279684 6194 280062
rect 583520 272234 584960 272324
rect 579662 272174 584960 272234
rect 579662 271826 579722 272174
rect 583520 272084 584960 272174
rect 576748 271766 579722 271826
rect -960 267202 480 267292
rect -960 267142 3066 267202
rect -960 267052 480 267142
rect 3006 267066 3066 267142
rect 3006 267006 6164 267066
rect 583520 258906 584960 258996
rect 576748 258846 584960 258906
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 6134 254146 6194 254388
rect -960 254086 6194 254146
rect -960 253996 480 254086
rect 576748 245926 579538 245986
rect 579478 245714 579538 245926
rect 579478 245654 579722 245714
rect 579662 245578 579722 245654
rect 583520 245578 584960 245668
rect 579662 245518 584960 245578
rect 583520 245428 584960 245518
rect 6134 241634 6194 241740
rect 3006 241574 6194 241634
rect -960 241090 480 241180
rect 3006 241090 3066 241574
rect -960 241030 3066 241090
rect -960 240940 480 241030
rect 576748 233006 583586 233066
rect 583526 232522 583586 233006
rect 583342 232476 583586 232522
rect 583342 232462 584960 232476
rect 583342 232386 583402 232462
rect 583520 232386 584960 232462
rect 583342 232326 584960 232386
rect 583520 232236 584960 232326
rect 3049 229122 3115 229125
rect 3049 229120 6164 229122
rect 3049 229064 3054 229120
rect 3110 229064 6164 229120
rect 3049 229062 6164 229064
rect 3049 229059 3115 229062
rect -960 228034 480 228124
rect 3049 228034 3115 228037
rect -960 228032 3115 228034
rect -960 227976 3054 228032
rect 3110 227976 3115 228032
rect -960 227974 3115 227976
rect -960 227884 480 227974
rect 3049 227971 3115 227974
rect 578509 220146 578575 220149
rect 576748 220144 578575 220146
rect 576748 220088 578514 220144
rect 578570 220088 578575 220144
rect 576748 220086 578575 220088
rect 578509 220083 578575 220086
rect 580901 219058 580967 219061
rect 583520 219058 584960 219148
rect 580901 219056 584960 219058
rect 580901 219000 580906 219056
rect 580962 219000 584960 219056
rect 580901 218998 584960 219000
rect 580901 218995 580967 218998
rect 583520 218908 584960 218998
rect 3049 216474 3115 216477
rect 3049 216472 6164 216474
rect 3049 216416 3054 216472
rect 3110 216416 6164 216472
rect 3049 216414 6164 216416
rect 3049 216411 3115 216414
rect -960 214978 480 215068
rect 3049 214978 3115 214981
rect -960 214976 3115 214978
rect -960 214920 3054 214976
rect 3110 214920 3115 214976
rect -960 214918 3115 214920
rect -960 214828 480 214918
rect 3049 214915 3115 214918
rect 579521 207226 579587 207229
rect 576748 207224 579587 207226
rect 576748 207168 579526 207224
rect 579582 207168 579587 207224
rect 576748 207166 579587 207168
rect 579521 207163 579587 207166
rect 579613 205730 579679 205733
rect 583520 205730 584960 205820
rect 579613 205728 584960 205730
rect 579613 205672 579618 205728
rect 579674 205672 584960 205728
rect 579613 205670 584960 205672
rect 579613 205667 579679 205670
rect 583520 205580 584960 205670
rect 3049 203826 3115 203829
rect 3049 203824 6164 203826
rect 3049 203768 3054 203824
rect 3110 203768 6164 203824
rect 3049 203766 6164 203768
rect 3049 203763 3115 203766
rect -960 201922 480 202012
rect 3049 201922 3115 201925
rect -960 201920 3115 201922
rect -960 201864 3054 201920
rect 3110 201864 3115 201920
rect -960 201862 3115 201864
rect -960 201772 480 201862
rect 3049 201859 3115 201862
rect 579521 194306 579587 194309
rect 576748 194304 579587 194306
rect 576748 194248 579526 194304
rect 579582 194248 579587 194304
rect 576748 194246 579587 194248
rect 579521 194243 579587 194246
rect 579613 192538 579679 192541
rect 583520 192538 584960 192628
rect 579613 192536 584960 192538
rect 579613 192480 579618 192536
rect 579674 192480 584960 192536
rect 579613 192478 584960 192480
rect 579613 192475 579679 192478
rect 583520 192388 584960 192478
rect 2957 191178 3023 191181
rect 2957 191176 6164 191178
rect 2957 191120 2962 191176
rect 3018 191120 6164 191176
rect 2957 191118 6164 191120
rect 2957 191115 3023 191118
rect -960 188866 480 188956
rect 2957 188866 3023 188869
rect -960 188864 3023 188866
rect -960 188808 2962 188864
rect 3018 188808 3023 188864
rect -960 188806 3023 188808
rect -960 188716 480 188806
rect 2957 188803 3023 188806
rect 578325 181386 578391 181389
rect 576748 181384 578391 181386
rect 576748 181328 578330 181384
rect 578386 181328 578391 181384
rect 576748 181326 578391 181328
rect 578325 181323 578391 181326
rect 580533 179210 580599 179213
rect 583520 179210 584960 179300
rect 580533 179208 584960 179210
rect 580533 179152 580538 179208
rect 580594 179152 584960 179208
rect 580533 179150 584960 179152
rect 580533 179147 580599 179150
rect 583520 179060 584960 179150
rect 2957 178530 3023 178533
rect 2957 178528 6164 178530
rect 2957 178472 2962 178528
rect 3018 178472 6164 178528
rect 2957 178470 6164 178472
rect 2957 178467 3023 178470
rect -960 175946 480 176036
rect 2957 175946 3023 175949
rect -960 175944 3023 175946
rect -960 175888 2962 175944
rect 3018 175888 3023 175944
rect -960 175886 3023 175888
rect -960 175796 480 175886
rect 2957 175883 3023 175886
rect 579521 168466 579587 168469
rect 576748 168464 579587 168466
rect 576748 168408 579526 168464
rect 579582 168408 579587 168464
rect 576748 168406 579587 168408
rect 579521 168403 579587 168406
rect 3049 165882 3115 165885
rect 579613 165882 579679 165885
rect 583520 165882 584960 165972
rect 3049 165880 6164 165882
rect 3049 165824 3054 165880
rect 3110 165824 6164 165880
rect 3049 165822 6164 165824
rect 579613 165880 584960 165882
rect 579613 165824 579618 165880
rect 579674 165824 584960 165880
rect 579613 165822 584960 165824
rect 3049 165819 3115 165822
rect 579613 165819 579679 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3049 162890 3115 162893
rect -960 162888 3115 162890
rect -960 162832 3054 162888
rect 3110 162832 3115 162888
rect -960 162830 3115 162832
rect -960 162740 480 162830
rect 3049 162827 3115 162830
rect 579521 155546 579587 155549
rect 576748 155544 579587 155546
rect 576748 155488 579526 155544
rect 579582 155488 579587 155544
rect 576748 155486 579587 155488
rect 579521 155483 579587 155486
rect 3049 153234 3115 153237
rect 3049 153232 6164 153234
rect 3049 153176 3054 153232
rect 3110 153176 6164 153232
rect 3049 153174 6164 153176
rect 3049 153171 3115 153174
rect 579613 152690 579679 152693
rect 583520 152690 584960 152780
rect 579613 152688 584960 152690
rect 579613 152632 579618 152688
rect 579674 152632 584960 152688
rect 579613 152630 584960 152632
rect 579613 152627 579679 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3049 149834 3115 149837
rect -960 149832 3115 149834
rect -960 149776 3054 149832
rect 3110 149776 3115 149832
rect -960 149774 3115 149776
rect -960 149684 480 149774
rect 3049 149771 3115 149774
rect 578785 142626 578851 142629
rect 576748 142624 578851 142626
rect 576748 142568 578790 142624
rect 578846 142568 578851 142624
rect 576748 142566 578851 142568
rect 578785 142563 578851 142566
rect 3049 140586 3115 140589
rect 3049 140584 6164 140586
rect 3049 140528 3054 140584
rect 3110 140528 6164 140584
rect 3049 140526 6164 140528
rect 3049 140523 3115 140526
rect 580717 139362 580783 139365
rect 583520 139362 584960 139452
rect 580717 139360 584960 139362
rect 580717 139304 580722 139360
rect 580778 139304 584960 139360
rect 580717 139302 584960 139304
rect 580717 139299 580783 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 3049 136778 3115 136781
rect -960 136776 3115 136778
rect -960 136720 3054 136776
rect 3110 136720 3115 136776
rect -960 136718 3115 136720
rect -960 136628 480 136718
rect 3049 136715 3115 136718
rect 579521 129706 579587 129709
rect 576748 129704 579587 129706
rect 576748 129648 579526 129704
rect 579582 129648 579587 129704
rect 576748 129646 579587 129648
rect 579521 129643 579587 129646
rect 3049 127938 3115 127941
rect 3049 127936 6164 127938
rect 3049 127880 3054 127936
rect 3110 127880 6164 127936
rect 3049 127878 6164 127880
rect 3049 127875 3115 127878
rect 579613 126034 579679 126037
rect 583520 126034 584960 126124
rect 579613 126032 584960 126034
rect 579613 125976 579618 126032
rect 579674 125976 584960 126032
rect 579613 125974 584960 125976
rect 579613 125971 579679 125974
rect 583520 125884 584960 125974
rect -960 123722 480 123812
rect 3049 123722 3115 123725
rect -960 123720 3115 123722
rect -960 123664 3054 123720
rect 3110 123664 3115 123720
rect -960 123662 3115 123664
rect -960 123572 480 123662
rect 3049 123659 3115 123662
rect 578325 116786 578391 116789
rect 576748 116784 578391 116786
rect 576748 116728 578330 116784
rect 578386 116728 578391 116784
rect 576748 116726 578391 116728
rect 578325 116723 578391 116726
rect 2957 115290 3023 115293
rect 2957 115288 6164 115290
rect 2957 115232 2962 115288
rect 3018 115232 6164 115288
rect 2957 115230 6164 115232
rect 2957 115227 3023 115230
rect 580257 112842 580323 112845
rect 583520 112842 584960 112932
rect 580257 112840 584960 112842
rect 580257 112784 580262 112840
rect 580318 112784 584960 112840
rect 580257 112782 584960 112784
rect 580257 112779 580323 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 2957 110666 3023 110669
rect -960 110664 3023 110666
rect -960 110608 2962 110664
rect 3018 110608 3023 110664
rect -960 110606 3023 110608
rect -960 110516 480 110606
rect 2957 110603 3023 110606
rect 579521 103866 579587 103869
rect 576748 103864 579587 103866
rect 576748 103808 579526 103864
rect 579582 103808 579587 103864
rect 576748 103806 579587 103808
rect 579521 103803 579587 103806
rect 3049 102642 3115 102645
rect 3049 102640 6164 102642
rect 3049 102584 3054 102640
rect 3110 102584 6164 102640
rect 3049 102582 6164 102584
rect 3049 102579 3115 102582
rect 579797 99514 579863 99517
rect 583520 99514 584960 99604
rect 579797 99512 584960 99514
rect 579797 99456 579802 99512
rect 579858 99456 584960 99512
rect 579797 99454 584960 99456
rect 579797 99451 579863 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 3049 97610 3115 97613
rect -960 97608 3115 97610
rect -960 97552 3054 97608
rect 3110 97552 3115 97608
rect -960 97550 3115 97552
rect -960 97460 480 97550
rect 3049 97547 3115 97550
rect 579521 90946 579587 90949
rect 576748 90944 579587 90946
rect 576748 90888 579526 90944
rect 579582 90888 579587 90944
rect 576748 90886 579587 90888
rect 579521 90883 579587 90886
rect 3049 89994 3115 89997
rect 3049 89992 6164 89994
rect 3049 89936 3054 89992
rect 3110 89936 6164 89992
rect 3049 89934 6164 89936
rect 3049 89931 3115 89934
rect 579613 86186 579679 86189
rect 583520 86186 584960 86276
rect 579613 86184 584960 86186
rect 579613 86128 579618 86184
rect 579674 86128 584960 86184
rect 579613 86126 584960 86128
rect 579613 86123 579679 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3049 84690 3115 84693
rect -960 84688 3115 84690
rect -960 84632 3054 84688
rect 3110 84632 3115 84688
rect -960 84630 3115 84632
rect -960 84540 480 84630
rect 3049 84627 3115 84630
rect 578877 78026 578943 78029
rect 576748 78024 578943 78026
rect 576748 77968 578882 78024
rect 578938 77968 578943 78024
rect 576748 77966 578943 77968
rect 578877 77963 578943 77966
rect 3417 77346 3483 77349
rect 3417 77344 6164 77346
rect 3417 77288 3422 77344
rect 3478 77288 6164 77344
rect 3417 77286 6164 77288
rect 3417 77283 3483 77286
rect 578877 72994 578943 72997
rect 583520 72994 584960 73084
rect 578877 72992 584960 72994
rect 578877 72936 578882 72992
rect 578938 72936 584960 72992
rect 578877 72934 584960 72936
rect 578877 72931 578943 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 578233 65106 578299 65109
rect 576748 65104 578299 65106
rect 576748 65048 578238 65104
rect 578294 65048 578299 65104
rect 576748 65046 578299 65048
rect 578233 65043 578299 65046
rect 3049 64698 3115 64701
rect 3049 64696 6164 64698
rect 3049 64640 3054 64696
rect 3110 64640 6164 64696
rect 3049 64638 6164 64640
rect 3049 64635 3115 64638
rect 580809 59666 580875 59669
rect 583520 59666 584960 59756
rect 580809 59664 584960 59666
rect 580809 59608 580814 59664
rect 580870 59608 584960 59664
rect 580809 59606 584960 59608
rect 580809 59603 580875 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3049 58578 3115 58581
rect -960 58576 3115 58578
rect -960 58520 3054 58576
rect 3110 58520 3115 58576
rect -960 58518 3115 58520
rect -960 58428 480 58518
rect 3049 58515 3115 58518
rect 579521 52186 579587 52189
rect 576748 52184 579587 52186
rect 576748 52128 579526 52184
rect 579582 52128 579587 52184
rect 576748 52126 579587 52128
rect 579521 52123 579587 52126
rect 3417 52050 3483 52053
rect 3417 52048 6164 52050
rect 3417 51992 3422 52048
rect 3478 51992 6164 52048
rect 3417 51990 6164 51992
rect 3417 51987 3483 51990
rect 579521 46338 579587 46341
rect 583520 46338 584960 46428
rect 579521 46336 584960 46338
rect 579521 46280 579526 46336
rect 579582 46280 584960 46336
rect 579521 46278 584960 46280
rect 579521 46275 579587 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 3417 39402 3483 39405
rect 3417 39400 6164 39402
rect 3417 39344 3422 39400
rect 3478 39344 6164 39400
rect 3417 39342 6164 39344
rect 3417 39339 3483 39342
rect 578877 39266 578943 39269
rect 576748 39264 578943 39266
rect 576748 39208 578882 39264
rect 578938 39208 578943 39264
rect 576748 39206 578943 39208
rect 578877 39203 578943 39206
rect 578877 33146 578943 33149
rect 583520 33146 584960 33236
rect 578877 33144 584960 33146
rect 578877 33088 578882 33144
rect 578938 33088 584960 33144
rect 578877 33086 584960 33088
rect 578877 33083 578943 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3417 32466 3483 32469
rect -960 32464 3483 32466
rect -960 32408 3422 32464
rect 3478 32408 3483 32464
rect -960 32406 3483 32408
rect -960 32316 480 32406
rect 3417 32403 3483 32406
rect 2957 26754 3023 26757
rect 2957 26752 6164 26754
rect 2957 26696 2962 26752
rect 3018 26696 6164 26752
rect 2957 26694 6164 26696
rect 2957 26691 3023 26694
rect 578233 26346 578299 26349
rect 576748 26344 578299 26346
rect 576748 26288 578238 26344
rect 578294 26288 578299 26344
rect 576748 26286 578299 26288
rect 578233 26283 578299 26286
rect 580625 19818 580691 19821
rect 583520 19818 584960 19908
rect 580625 19816 584960 19818
rect 580625 19760 580630 19816
rect 580686 19760 584960 19816
rect 580625 19758 584960 19760
rect 580625 19755 580691 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 2957 19410 3023 19413
rect -960 19408 3023 19410
rect -960 19352 2962 19408
rect 3018 19352 3023 19408
rect -960 19350 3023 19352
rect -960 19260 480 19350
rect 2957 19347 3023 19350
rect 3417 14106 3483 14109
rect 3417 14104 6164 14106
rect 3417 14048 3422 14104
rect 3478 14048 6164 14104
rect 3417 14046 6164 14048
rect 3417 14043 3483 14046
rect 578877 13426 578943 13429
rect 576748 13424 578943 13426
rect 576748 13368 578882 13424
rect 578938 13368 578943 13424
rect 576748 13366 578943 13368
rect 578877 13363 578943 13366
rect 578877 6626 578943 6629
rect 583520 6626 584960 6716
rect 578877 6624 584960 6626
rect -960 6490 480 6580
rect 578877 6568 578882 6624
rect 578938 6568 584960 6624
rect 578877 6566 584960 6568
rect 578877 6563 578943 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 539133 3770 539199 3773
rect 557349 3770 557415 3773
rect 539133 3768 557415 3770
rect 539133 3712 539138 3768
rect 539194 3712 557354 3768
rect 557410 3712 557415 3768
rect 539133 3710 557415 3712
rect 539133 3707 539199 3710
rect 557349 3707 557415 3710
rect 552381 3634 552447 3637
rect 571517 3634 571583 3637
rect 552381 3632 571583 3634
rect 552381 3576 552386 3632
rect 552442 3576 571522 3632
rect 571578 3576 571583 3632
rect 552381 3574 571583 3576
rect 552381 3571 552447 3574
rect 571517 3571 571583 3574
rect 20621 3498 20687 3501
rect 37917 3498 37983 3501
rect 20621 3496 37983 3498
rect 20621 3440 20626 3496
rect 20682 3440 37922 3496
rect 37978 3440 37983 3496
rect 20621 3438 37983 3440
rect 20621 3435 20687 3438
rect 37917 3435 37983 3438
rect 521469 3498 521535 3501
rect 538397 3498 538463 3501
rect 521469 3496 538463 3498
rect 521469 3440 521474 3496
rect 521530 3440 538402 3496
rect 538458 3440 538463 3496
rect 521469 3438 538463 3440
rect 521469 3435 521535 3438
rect 538397 3435 538463 3438
rect 555693 3498 555759 3501
rect 575105 3498 575171 3501
rect 555693 3496 575171 3498
rect 555693 3440 555698 3496
rect 555754 3440 575110 3496
rect 575166 3440 575171 3496
rect 555693 3438 575171 3440
rect 555693 3435 555759 3438
rect 575105 3435 575171 3438
rect 5257 3362 5323 3365
rect 23565 3362 23631 3365
rect 5257 3360 23631 3362
rect 5257 3304 5262 3360
rect 5318 3304 23570 3360
rect 23626 3304 23631 3360
rect 5257 3302 23631 3304
rect 5257 3299 5323 3302
rect 23565 3299 23631 3302
rect 28901 3362 28967 3365
rect 45645 3362 45711 3365
rect 28901 3360 45711 3362
rect 28901 3304 28906 3360
rect 28962 3304 45650 3360
rect 45706 3304 45711 3360
rect 28901 3302 45711 3304
rect 28901 3299 28967 3302
rect 45645 3299 45711 3302
rect 538029 3362 538095 3365
rect 556153 3362 556219 3365
rect 538029 3360 556219 3362
rect 538029 3304 538034 3360
rect 538090 3304 556158 3360
rect 556214 3304 556219 3360
rect 538029 3302 556219 3304
rect 538029 3299 538095 3302
rect 556153 3299 556219 3302
rect 560109 3362 560175 3365
rect 579797 3362 579863 3365
rect 560109 3360 579863 3362
rect 560109 3304 560114 3360
rect 560170 3304 579802 3360
rect 579858 3304 579863 3360
rect 560109 3302 579863 3304
rect 560109 3299 560175 3302
rect 579797 3299 579863 3302
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 677494 -8106 711002
rect -8726 677258 -8694 677494
rect -8458 677258 -8374 677494
rect -8138 677258 -8106 677494
rect -8726 677174 -8106 677258
rect -8726 676938 -8694 677174
rect -8458 676938 -8374 677174
rect -8138 676938 -8106 677174
rect -8726 641494 -8106 676938
rect -8726 641258 -8694 641494
rect -8458 641258 -8374 641494
rect -8138 641258 -8106 641494
rect -8726 641174 -8106 641258
rect -8726 640938 -8694 641174
rect -8458 640938 -8374 641174
rect -8138 640938 -8106 641174
rect -8726 605494 -8106 640938
rect -8726 605258 -8694 605494
rect -8458 605258 -8374 605494
rect -8138 605258 -8106 605494
rect -8726 605174 -8106 605258
rect -8726 604938 -8694 605174
rect -8458 604938 -8374 605174
rect -8138 604938 -8106 605174
rect -8726 569494 -8106 604938
rect -8726 569258 -8694 569494
rect -8458 569258 -8374 569494
rect -8138 569258 -8106 569494
rect -8726 569174 -8106 569258
rect -8726 568938 -8694 569174
rect -8458 568938 -8374 569174
rect -8138 568938 -8106 569174
rect -8726 533494 -8106 568938
rect -8726 533258 -8694 533494
rect -8458 533258 -8374 533494
rect -8138 533258 -8106 533494
rect -8726 533174 -8106 533258
rect -8726 532938 -8694 533174
rect -8458 532938 -8374 533174
rect -8138 532938 -8106 533174
rect -8726 497494 -8106 532938
rect -8726 497258 -8694 497494
rect -8458 497258 -8374 497494
rect -8138 497258 -8106 497494
rect -8726 497174 -8106 497258
rect -8726 496938 -8694 497174
rect -8458 496938 -8374 497174
rect -8138 496938 -8106 497174
rect -8726 461494 -8106 496938
rect -8726 461258 -8694 461494
rect -8458 461258 -8374 461494
rect -8138 461258 -8106 461494
rect -8726 461174 -8106 461258
rect -8726 460938 -8694 461174
rect -8458 460938 -8374 461174
rect -8138 460938 -8106 461174
rect -8726 425494 -8106 460938
rect -8726 425258 -8694 425494
rect -8458 425258 -8374 425494
rect -8138 425258 -8106 425494
rect -8726 425174 -8106 425258
rect -8726 424938 -8694 425174
rect -8458 424938 -8374 425174
rect -8138 424938 -8106 425174
rect -8726 389494 -8106 424938
rect -8726 389258 -8694 389494
rect -8458 389258 -8374 389494
rect -8138 389258 -8106 389494
rect -8726 389174 -8106 389258
rect -8726 388938 -8694 389174
rect -8458 388938 -8374 389174
rect -8138 388938 -8106 389174
rect -8726 353494 -8106 388938
rect -8726 353258 -8694 353494
rect -8458 353258 -8374 353494
rect -8138 353258 -8106 353494
rect -8726 353174 -8106 353258
rect -8726 352938 -8694 353174
rect -8458 352938 -8374 353174
rect -8138 352938 -8106 353174
rect -8726 317494 -8106 352938
rect -8726 317258 -8694 317494
rect -8458 317258 -8374 317494
rect -8138 317258 -8106 317494
rect -8726 317174 -8106 317258
rect -8726 316938 -8694 317174
rect -8458 316938 -8374 317174
rect -8138 316938 -8106 317174
rect -8726 281494 -8106 316938
rect -8726 281258 -8694 281494
rect -8458 281258 -8374 281494
rect -8138 281258 -8106 281494
rect -8726 281174 -8106 281258
rect -8726 280938 -8694 281174
rect -8458 280938 -8374 281174
rect -8138 280938 -8106 281174
rect -8726 245494 -8106 280938
rect -8726 245258 -8694 245494
rect -8458 245258 -8374 245494
rect -8138 245258 -8106 245494
rect -8726 245174 -8106 245258
rect -8726 244938 -8694 245174
rect -8458 244938 -8374 245174
rect -8138 244938 -8106 245174
rect -8726 209494 -8106 244938
rect -8726 209258 -8694 209494
rect -8458 209258 -8374 209494
rect -8138 209258 -8106 209494
rect -8726 209174 -8106 209258
rect -8726 208938 -8694 209174
rect -8458 208938 -8374 209174
rect -8138 208938 -8106 209174
rect -8726 173494 -8106 208938
rect -8726 173258 -8694 173494
rect -8458 173258 -8374 173494
rect -8138 173258 -8106 173494
rect -8726 173174 -8106 173258
rect -8726 172938 -8694 173174
rect -8458 172938 -8374 173174
rect -8138 172938 -8106 173174
rect -8726 137494 -8106 172938
rect -8726 137258 -8694 137494
rect -8458 137258 -8374 137494
rect -8138 137258 -8106 137494
rect -8726 137174 -8106 137258
rect -8726 136938 -8694 137174
rect -8458 136938 -8374 137174
rect -8138 136938 -8106 137174
rect -8726 101494 -8106 136938
rect -8726 101258 -8694 101494
rect -8458 101258 -8374 101494
rect -8138 101258 -8106 101494
rect -8726 101174 -8106 101258
rect -8726 100938 -8694 101174
rect -8458 100938 -8374 101174
rect -8138 100938 -8106 101174
rect -8726 65494 -8106 100938
rect -8726 65258 -8694 65494
rect -8458 65258 -8374 65494
rect -8138 65258 -8106 65494
rect -8726 65174 -8106 65258
rect -8726 64938 -8694 65174
rect -8458 64938 -8374 65174
rect -8138 64938 -8106 65174
rect -8726 29494 -8106 64938
rect -8726 29258 -8694 29494
rect -8458 29258 -8374 29494
rect -8138 29258 -8106 29494
rect -8726 29174 -8106 29258
rect -8726 28938 -8694 29174
rect -8458 28938 -8374 29174
rect -8138 28938 -8106 29174
rect -8726 -7066 -8106 28938
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 673774 -7146 710042
rect -7766 673538 -7734 673774
rect -7498 673538 -7414 673774
rect -7178 673538 -7146 673774
rect -7766 673454 -7146 673538
rect -7766 673218 -7734 673454
rect -7498 673218 -7414 673454
rect -7178 673218 -7146 673454
rect -7766 637774 -7146 673218
rect -7766 637538 -7734 637774
rect -7498 637538 -7414 637774
rect -7178 637538 -7146 637774
rect -7766 637454 -7146 637538
rect -7766 637218 -7734 637454
rect -7498 637218 -7414 637454
rect -7178 637218 -7146 637454
rect -7766 601774 -7146 637218
rect -7766 601538 -7734 601774
rect -7498 601538 -7414 601774
rect -7178 601538 -7146 601774
rect -7766 601454 -7146 601538
rect -7766 601218 -7734 601454
rect -7498 601218 -7414 601454
rect -7178 601218 -7146 601454
rect -7766 565774 -7146 601218
rect -7766 565538 -7734 565774
rect -7498 565538 -7414 565774
rect -7178 565538 -7146 565774
rect -7766 565454 -7146 565538
rect -7766 565218 -7734 565454
rect -7498 565218 -7414 565454
rect -7178 565218 -7146 565454
rect -7766 529774 -7146 565218
rect -7766 529538 -7734 529774
rect -7498 529538 -7414 529774
rect -7178 529538 -7146 529774
rect -7766 529454 -7146 529538
rect -7766 529218 -7734 529454
rect -7498 529218 -7414 529454
rect -7178 529218 -7146 529454
rect -7766 493774 -7146 529218
rect -7766 493538 -7734 493774
rect -7498 493538 -7414 493774
rect -7178 493538 -7146 493774
rect -7766 493454 -7146 493538
rect -7766 493218 -7734 493454
rect -7498 493218 -7414 493454
rect -7178 493218 -7146 493454
rect -7766 457774 -7146 493218
rect -7766 457538 -7734 457774
rect -7498 457538 -7414 457774
rect -7178 457538 -7146 457774
rect -7766 457454 -7146 457538
rect -7766 457218 -7734 457454
rect -7498 457218 -7414 457454
rect -7178 457218 -7146 457454
rect -7766 421774 -7146 457218
rect -7766 421538 -7734 421774
rect -7498 421538 -7414 421774
rect -7178 421538 -7146 421774
rect -7766 421454 -7146 421538
rect -7766 421218 -7734 421454
rect -7498 421218 -7414 421454
rect -7178 421218 -7146 421454
rect -7766 385774 -7146 421218
rect -7766 385538 -7734 385774
rect -7498 385538 -7414 385774
rect -7178 385538 -7146 385774
rect -7766 385454 -7146 385538
rect -7766 385218 -7734 385454
rect -7498 385218 -7414 385454
rect -7178 385218 -7146 385454
rect -7766 349774 -7146 385218
rect -7766 349538 -7734 349774
rect -7498 349538 -7414 349774
rect -7178 349538 -7146 349774
rect -7766 349454 -7146 349538
rect -7766 349218 -7734 349454
rect -7498 349218 -7414 349454
rect -7178 349218 -7146 349454
rect -7766 313774 -7146 349218
rect -7766 313538 -7734 313774
rect -7498 313538 -7414 313774
rect -7178 313538 -7146 313774
rect -7766 313454 -7146 313538
rect -7766 313218 -7734 313454
rect -7498 313218 -7414 313454
rect -7178 313218 -7146 313454
rect -7766 277774 -7146 313218
rect -7766 277538 -7734 277774
rect -7498 277538 -7414 277774
rect -7178 277538 -7146 277774
rect -7766 277454 -7146 277538
rect -7766 277218 -7734 277454
rect -7498 277218 -7414 277454
rect -7178 277218 -7146 277454
rect -7766 241774 -7146 277218
rect -7766 241538 -7734 241774
rect -7498 241538 -7414 241774
rect -7178 241538 -7146 241774
rect -7766 241454 -7146 241538
rect -7766 241218 -7734 241454
rect -7498 241218 -7414 241454
rect -7178 241218 -7146 241454
rect -7766 205774 -7146 241218
rect -7766 205538 -7734 205774
rect -7498 205538 -7414 205774
rect -7178 205538 -7146 205774
rect -7766 205454 -7146 205538
rect -7766 205218 -7734 205454
rect -7498 205218 -7414 205454
rect -7178 205218 -7146 205454
rect -7766 169774 -7146 205218
rect -7766 169538 -7734 169774
rect -7498 169538 -7414 169774
rect -7178 169538 -7146 169774
rect -7766 169454 -7146 169538
rect -7766 169218 -7734 169454
rect -7498 169218 -7414 169454
rect -7178 169218 -7146 169454
rect -7766 133774 -7146 169218
rect -7766 133538 -7734 133774
rect -7498 133538 -7414 133774
rect -7178 133538 -7146 133774
rect -7766 133454 -7146 133538
rect -7766 133218 -7734 133454
rect -7498 133218 -7414 133454
rect -7178 133218 -7146 133454
rect -7766 97774 -7146 133218
rect -7766 97538 -7734 97774
rect -7498 97538 -7414 97774
rect -7178 97538 -7146 97774
rect -7766 97454 -7146 97538
rect -7766 97218 -7734 97454
rect -7498 97218 -7414 97454
rect -7178 97218 -7146 97454
rect -7766 61774 -7146 97218
rect -7766 61538 -7734 61774
rect -7498 61538 -7414 61774
rect -7178 61538 -7146 61774
rect -7766 61454 -7146 61538
rect -7766 61218 -7734 61454
rect -7498 61218 -7414 61454
rect -7178 61218 -7146 61454
rect -7766 25774 -7146 61218
rect -7766 25538 -7734 25774
rect -7498 25538 -7414 25774
rect -7178 25538 -7146 25774
rect -7766 25454 -7146 25538
rect -7766 25218 -7734 25454
rect -7498 25218 -7414 25454
rect -7178 25218 -7146 25454
rect -7766 -6106 -7146 25218
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 670054 -6186 709082
rect -6806 669818 -6774 670054
rect -6538 669818 -6454 670054
rect -6218 669818 -6186 670054
rect -6806 669734 -6186 669818
rect -6806 669498 -6774 669734
rect -6538 669498 -6454 669734
rect -6218 669498 -6186 669734
rect -6806 634054 -6186 669498
rect -6806 633818 -6774 634054
rect -6538 633818 -6454 634054
rect -6218 633818 -6186 634054
rect -6806 633734 -6186 633818
rect -6806 633498 -6774 633734
rect -6538 633498 -6454 633734
rect -6218 633498 -6186 633734
rect -6806 598054 -6186 633498
rect -6806 597818 -6774 598054
rect -6538 597818 -6454 598054
rect -6218 597818 -6186 598054
rect -6806 597734 -6186 597818
rect -6806 597498 -6774 597734
rect -6538 597498 -6454 597734
rect -6218 597498 -6186 597734
rect -6806 562054 -6186 597498
rect -6806 561818 -6774 562054
rect -6538 561818 -6454 562054
rect -6218 561818 -6186 562054
rect -6806 561734 -6186 561818
rect -6806 561498 -6774 561734
rect -6538 561498 -6454 561734
rect -6218 561498 -6186 561734
rect -6806 526054 -6186 561498
rect -6806 525818 -6774 526054
rect -6538 525818 -6454 526054
rect -6218 525818 -6186 526054
rect -6806 525734 -6186 525818
rect -6806 525498 -6774 525734
rect -6538 525498 -6454 525734
rect -6218 525498 -6186 525734
rect -6806 490054 -6186 525498
rect -6806 489818 -6774 490054
rect -6538 489818 -6454 490054
rect -6218 489818 -6186 490054
rect -6806 489734 -6186 489818
rect -6806 489498 -6774 489734
rect -6538 489498 -6454 489734
rect -6218 489498 -6186 489734
rect -6806 454054 -6186 489498
rect -6806 453818 -6774 454054
rect -6538 453818 -6454 454054
rect -6218 453818 -6186 454054
rect -6806 453734 -6186 453818
rect -6806 453498 -6774 453734
rect -6538 453498 -6454 453734
rect -6218 453498 -6186 453734
rect -6806 418054 -6186 453498
rect -6806 417818 -6774 418054
rect -6538 417818 -6454 418054
rect -6218 417818 -6186 418054
rect -6806 417734 -6186 417818
rect -6806 417498 -6774 417734
rect -6538 417498 -6454 417734
rect -6218 417498 -6186 417734
rect -6806 382054 -6186 417498
rect -6806 381818 -6774 382054
rect -6538 381818 -6454 382054
rect -6218 381818 -6186 382054
rect -6806 381734 -6186 381818
rect -6806 381498 -6774 381734
rect -6538 381498 -6454 381734
rect -6218 381498 -6186 381734
rect -6806 346054 -6186 381498
rect -6806 345818 -6774 346054
rect -6538 345818 -6454 346054
rect -6218 345818 -6186 346054
rect -6806 345734 -6186 345818
rect -6806 345498 -6774 345734
rect -6538 345498 -6454 345734
rect -6218 345498 -6186 345734
rect -6806 310054 -6186 345498
rect -6806 309818 -6774 310054
rect -6538 309818 -6454 310054
rect -6218 309818 -6186 310054
rect -6806 309734 -6186 309818
rect -6806 309498 -6774 309734
rect -6538 309498 -6454 309734
rect -6218 309498 -6186 309734
rect -6806 274054 -6186 309498
rect -6806 273818 -6774 274054
rect -6538 273818 -6454 274054
rect -6218 273818 -6186 274054
rect -6806 273734 -6186 273818
rect -6806 273498 -6774 273734
rect -6538 273498 -6454 273734
rect -6218 273498 -6186 273734
rect -6806 238054 -6186 273498
rect -6806 237818 -6774 238054
rect -6538 237818 -6454 238054
rect -6218 237818 -6186 238054
rect -6806 237734 -6186 237818
rect -6806 237498 -6774 237734
rect -6538 237498 -6454 237734
rect -6218 237498 -6186 237734
rect -6806 202054 -6186 237498
rect -6806 201818 -6774 202054
rect -6538 201818 -6454 202054
rect -6218 201818 -6186 202054
rect -6806 201734 -6186 201818
rect -6806 201498 -6774 201734
rect -6538 201498 -6454 201734
rect -6218 201498 -6186 201734
rect -6806 166054 -6186 201498
rect -6806 165818 -6774 166054
rect -6538 165818 -6454 166054
rect -6218 165818 -6186 166054
rect -6806 165734 -6186 165818
rect -6806 165498 -6774 165734
rect -6538 165498 -6454 165734
rect -6218 165498 -6186 165734
rect -6806 130054 -6186 165498
rect -6806 129818 -6774 130054
rect -6538 129818 -6454 130054
rect -6218 129818 -6186 130054
rect -6806 129734 -6186 129818
rect -6806 129498 -6774 129734
rect -6538 129498 -6454 129734
rect -6218 129498 -6186 129734
rect -6806 94054 -6186 129498
rect -6806 93818 -6774 94054
rect -6538 93818 -6454 94054
rect -6218 93818 -6186 94054
rect -6806 93734 -6186 93818
rect -6806 93498 -6774 93734
rect -6538 93498 -6454 93734
rect -6218 93498 -6186 93734
rect -6806 58054 -6186 93498
rect -6806 57818 -6774 58054
rect -6538 57818 -6454 58054
rect -6218 57818 -6186 58054
rect -6806 57734 -6186 57818
rect -6806 57498 -6774 57734
rect -6538 57498 -6454 57734
rect -6218 57498 -6186 57734
rect -6806 22054 -6186 57498
rect -6806 21818 -6774 22054
rect -6538 21818 -6454 22054
rect -6218 21818 -6186 22054
rect -6806 21734 -6186 21818
rect -6806 21498 -6774 21734
rect -6538 21498 -6454 21734
rect -6218 21498 -6186 21734
rect -6806 -5146 -6186 21498
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 666334 -5226 708122
rect -5846 666098 -5814 666334
rect -5578 666098 -5494 666334
rect -5258 666098 -5226 666334
rect -5846 666014 -5226 666098
rect -5846 665778 -5814 666014
rect -5578 665778 -5494 666014
rect -5258 665778 -5226 666014
rect -5846 630334 -5226 665778
rect -5846 630098 -5814 630334
rect -5578 630098 -5494 630334
rect -5258 630098 -5226 630334
rect -5846 630014 -5226 630098
rect -5846 629778 -5814 630014
rect -5578 629778 -5494 630014
rect -5258 629778 -5226 630014
rect -5846 594334 -5226 629778
rect -5846 594098 -5814 594334
rect -5578 594098 -5494 594334
rect -5258 594098 -5226 594334
rect -5846 594014 -5226 594098
rect -5846 593778 -5814 594014
rect -5578 593778 -5494 594014
rect -5258 593778 -5226 594014
rect -5846 558334 -5226 593778
rect -5846 558098 -5814 558334
rect -5578 558098 -5494 558334
rect -5258 558098 -5226 558334
rect -5846 558014 -5226 558098
rect -5846 557778 -5814 558014
rect -5578 557778 -5494 558014
rect -5258 557778 -5226 558014
rect -5846 522334 -5226 557778
rect -5846 522098 -5814 522334
rect -5578 522098 -5494 522334
rect -5258 522098 -5226 522334
rect -5846 522014 -5226 522098
rect -5846 521778 -5814 522014
rect -5578 521778 -5494 522014
rect -5258 521778 -5226 522014
rect -5846 486334 -5226 521778
rect -5846 486098 -5814 486334
rect -5578 486098 -5494 486334
rect -5258 486098 -5226 486334
rect -5846 486014 -5226 486098
rect -5846 485778 -5814 486014
rect -5578 485778 -5494 486014
rect -5258 485778 -5226 486014
rect -5846 450334 -5226 485778
rect -5846 450098 -5814 450334
rect -5578 450098 -5494 450334
rect -5258 450098 -5226 450334
rect -5846 450014 -5226 450098
rect -5846 449778 -5814 450014
rect -5578 449778 -5494 450014
rect -5258 449778 -5226 450014
rect -5846 414334 -5226 449778
rect -5846 414098 -5814 414334
rect -5578 414098 -5494 414334
rect -5258 414098 -5226 414334
rect -5846 414014 -5226 414098
rect -5846 413778 -5814 414014
rect -5578 413778 -5494 414014
rect -5258 413778 -5226 414014
rect -5846 378334 -5226 413778
rect -5846 378098 -5814 378334
rect -5578 378098 -5494 378334
rect -5258 378098 -5226 378334
rect -5846 378014 -5226 378098
rect -5846 377778 -5814 378014
rect -5578 377778 -5494 378014
rect -5258 377778 -5226 378014
rect -5846 342334 -5226 377778
rect -5846 342098 -5814 342334
rect -5578 342098 -5494 342334
rect -5258 342098 -5226 342334
rect -5846 342014 -5226 342098
rect -5846 341778 -5814 342014
rect -5578 341778 -5494 342014
rect -5258 341778 -5226 342014
rect -5846 306334 -5226 341778
rect -5846 306098 -5814 306334
rect -5578 306098 -5494 306334
rect -5258 306098 -5226 306334
rect -5846 306014 -5226 306098
rect -5846 305778 -5814 306014
rect -5578 305778 -5494 306014
rect -5258 305778 -5226 306014
rect -5846 270334 -5226 305778
rect -5846 270098 -5814 270334
rect -5578 270098 -5494 270334
rect -5258 270098 -5226 270334
rect -5846 270014 -5226 270098
rect -5846 269778 -5814 270014
rect -5578 269778 -5494 270014
rect -5258 269778 -5226 270014
rect -5846 234334 -5226 269778
rect -5846 234098 -5814 234334
rect -5578 234098 -5494 234334
rect -5258 234098 -5226 234334
rect -5846 234014 -5226 234098
rect -5846 233778 -5814 234014
rect -5578 233778 -5494 234014
rect -5258 233778 -5226 234014
rect -5846 198334 -5226 233778
rect -5846 198098 -5814 198334
rect -5578 198098 -5494 198334
rect -5258 198098 -5226 198334
rect -5846 198014 -5226 198098
rect -5846 197778 -5814 198014
rect -5578 197778 -5494 198014
rect -5258 197778 -5226 198014
rect -5846 162334 -5226 197778
rect -5846 162098 -5814 162334
rect -5578 162098 -5494 162334
rect -5258 162098 -5226 162334
rect -5846 162014 -5226 162098
rect -5846 161778 -5814 162014
rect -5578 161778 -5494 162014
rect -5258 161778 -5226 162014
rect -5846 126334 -5226 161778
rect -5846 126098 -5814 126334
rect -5578 126098 -5494 126334
rect -5258 126098 -5226 126334
rect -5846 126014 -5226 126098
rect -5846 125778 -5814 126014
rect -5578 125778 -5494 126014
rect -5258 125778 -5226 126014
rect -5846 90334 -5226 125778
rect -5846 90098 -5814 90334
rect -5578 90098 -5494 90334
rect -5258 90098 -5226 90334
rect -5846 90014 -5226 90098
rect -5846 89778 -5814 90014
rect -5578 89778 -5494 90014
rect -5258 89778 -5226 90014
rect -5846 54334 -5226 89778
rect -5846 54098 -5814 54334
rect -5578 54098 -5494 54334
rect -5258 54098 -5226 54334
rect -5846 54014 -5226 54098
rect -5846 53778 -5814 54014
rect -5578 53778 -5494 54014
rect -5258 53778 -5226 54014
rect -5846 18334 -5226 53778
rect -5846 18098 -5814 18334
rect -5578 18098 -5494 18334
rect -5258 18098 -5226 18334
rect -5846 18014 -5226 18098
rect -5846 17778 -5814 18014
rect -5578 17778 -5494 18014
rect -5258 17778 -5226 18014
rect -5846 -4186 -5226 17778
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 698614 -4266 707162
rect -4886 698378 -4854 698614
rect -4618 698378 -4534 698614
rect -4298 698378 -4266 698614
rect -4886 698294 -4266 698378
rect -4886 698058 -4854 698294
rect -4618 698058 -4534 698294
rect -4298 698058 -4266 698294
rect -4886 662614 -4266 698058
rect -4886 662378 -4854 662614
rect -4618 662378 -4534 662614
rect -4298 662378 -4266 662614
rect -4886 662294 -4266 662378
rect -4886 662058 -4854 662294
rect -4618 662058 -4534 662294
rect -4298 662058 -4266 662294
rect -4886 626614 -4266 662058
rect -4886 626378 -4854 626614
rect -4618 626378 -4534 626614
rect -4298 626378 -4266 626614
rect -4886 626294 -4266 626378
rect -4886 626058 -4854 626294
rect -4618 626058 -4534 626294
rect -4298 626058 -4266 626294
rect -4886 590614 -4266 626058
rect -4886 590378 -4854 590614
rect -4618 590378 -4534 590614
rect -4298 590378 -4266 590614
rect -4886 590294 -4266 590378
rect -4886 590058 -4854 590294
rect -4618 590058 -4534 590294
rect -4298 590058 -4266 590294
rect -4886 554614 -4266 590058
rect -4886 554378 -4854 554614
rect -4618 554378 -4534 554614
rect -4298 554378 -4266 554614
rect -4886 554294 -4266 554378
rect -4886 554058 -4854 554294
rect -4618 554058 -4534 554294
rect -4298 554058 -4266 554294
rect -4886 518614 -4266 554058
rect -4886 518378 -4854 518614
rect -4618 518378 -4534 518614
rect -4298 518378 -4266 518614
rect -4886 518294 -4266 518378
rect -4886 518058 -4854 518294
rect -4618 518058 -4534 518294
rect -4298 518058 -4266 518294
rect -4886 482614 -4266 518058
rect -4886 482378 -4854 482614
rect -4618 482378 -4534 482614
rect -4298 482378 -4266 482614
rect -4886 482294 -4266 482378
rect -4886 482058 -4854 482294
rect -4618 482058 -4534 482294
rect -4298 482058 -4266 482294
rect -4886 446614 -4266 482058
rect -4886 446378 -4854 446614
rect -4618 446378 -4534 446614
rect -4298 446378 -4266 446614
rect -4886 446294 -4266 446378
rect -4886 446058 -4854 446294
rect -4618 446058 -4534 446294
rect -4298 446058 -4266 446294
rect -4886 410614 -4266 446058
rect -4886 410378 -4854 410614
rect -4618 410378 -4534 410614
rect -4298 410378 -4266 410614
rect -4886 410294 -4266 410378
rect -4886 410058 -4854 410294
rect -4618 410058 -4534 410294
rect -4298 410058 -4266 410294
rect -4886 374614 -4266 410058
rect -4886 374378 -4854 374614
rect -4618 374378 -4534 374614
rect -4298 374378 -4266 374614
rect -4886 374294 -4266 374378
rect -4886 374058 -4854 374294
rect -4618 374058 -4534 374294
rect -4298 374058 -4266 374294
rect -4886 338614 -4266 374058
rect -4886 338378 -4854 338614
rect -4618 338378 -4534 338614
rect -4298 338378 -4266 338614
rect -4886 338294 -4266 338378
rect -4886 338058 -4854 338294
rect -4618 338058 -4534 338294
rect -4298 338058 -4266 338294
rect -4886 302614 -4266 338058
rect -4886 302378 -4854 302614
rect -4618 302378 -4534 302614
rect -4298 302378 -4266 302614
rect -4886 302294 -4266 302378
rect -4886 302058 -4854 302294
rect -4618 302058 -4534 302294
rect -4298 302058 -4266 302294
rect -4886 266614 -4266 302058
rect -4886 266378 -4854 266614
rect -4618 266378 -4534 266614
rect -4298 266378 -4266 266614
rect -4886 266294 -4266 266378
rect -4886 266058 -4854 266294
rect -4618 266058 -4534 266294
rect -4298 266058 -4266 266294
rect -4886 230614 -4266 266058
rect -4886 230378 -4854 230614
rect -4618 230378 -4534 230614
rect -4298 230378 -4266 230614
rect -4886 230294 -4266 230378
rect -4886 230058 -4854 230294
rect -4618 230058 -4534 230294
rect -4298 230058 -4266 230294
rect -4886 194614 -4266 230058
rect -4886 194378 -4854 194614
rect -4618 194378 -4534 194614
rect -4298 194378 -4266 194614
rect -4886 194294 -4266 194378
rect -4886 194058 -4854 194294
rect -4618 194058 -4534 194294
rect -4298 194058 -4266 194294
rect -4886 158614 -4266 194058
rect -4886 158378 -4854 158614
rect -4618 158378 -4534 158614
rect -4298 158378 -4266 158614
rect -4886 158294 -4266 158378
rect -4886 158058 -4854 158294
rect -4618 158058 -4534 158294
rect -4298 158058 -4266 158294
rect -4886 122614 -4266 158058
rect -4886 122378 -4854 122614
rect -4618 122378 -4534 122614
rect -4298 122378 -4266 122614
rect -4886 122294 -4266 122378
rect -4886 122058 -4854 122294
rect -4618 122058 -4534 122294
rect -4298 122058 -4266 122294
rect -4886 86614 -4266 122058
rect -4886 86378 -4854 86614
rect -4618 86378 -4534 86614
rect -4298 86378 -4266 86614
rect -4886 86294 -4266 86378
rect -4886 86058 -4854 86294
rect -4618 86058 -4534 86294
rect -4298 86058 -4266 86294
rect -4886 50614 -4266 86058
rect -4886 50378 -4854 50614
rect -4618 50378 -4534 50614
rect -4298 50378 -4266 50614
rect -4886 50294 -4266 50378
rect -4886 50058 -4854 50294
rect -4618 50058 -4534 50294
rect -4298 50058 -4266 50294
rect -4886 14614 -4266 50058
rect -4886 14378 -4854 14614
rect -4618 14378 -4534 14614
rect -4298 14378 -4266 14614
rect -4886 14294 -4266 14378
rect -4886 14058 -4854 14294
rect -4618 14058 -4534 14294
rect -4298 14058 -4266 14294
rect -4886 -3226 -4266 14058
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 694894 -3306 706202
rect -3926 694658 -3894 694894
rect -3658 694658 -3574 694894
rect -3338 694658 -3306 694894
rect -3926 694574 -3306 694658
rect -3926 694338 -3894 694574
rect -3658 694338 -3574 694574
rect -3338 694338 -3306 694574
rect -3926 658894 -3306 694338
rect -3926 658658 -3894 658894
rect -3658 658658 -3574 658894
rect -3338 658658 -3306 658894
rect -3926 658574 -3306 658658
rect -3926 658338 -3894 658574
rect -3658 658338 -3574 658574
rect -3338 658338 -3306 658574
rect -3926 622894 -3306 658338
rect -3926 622658 -3894 622894
rect -3658 622658 -3574 622894
rect -3338 622658 -3306 622894
rect -3926 622574 -3306 622658
rect -3926 622338 -3894 622574
rect -3658 622338 -3574 622574
rect -3338 622338 -3306 622574
rect -3926 586894 -3306 622338
rect -3926 586658 -3894 586894
rect -3658 586658 -3574 586894
rect -3338 586658 -3306 586894
rect -3926 586574 -3306 586658
rect -3926 586338 -3894 586574
rect -3658 586338 -3574 586574
rect -3338 586338 -3306 586574
rect -3926 550894 -3306 586338
rect -3926 550658 -3894 550894
rect -3658 550658 -3574 550894
rect -3338 550658 -3306 550894
rect -3926 550574 -3306 550658
rect -3926 550338 -3894 550574
rect -3658 550338 -3574 550574
rect -3338 550338 -3306 550574
rect -3926 514894 -3306 550338
rect -3926 514658 -3894 514894
rect -3658 514658 -3574 514894
rect -3338 514658 -3306 514894
rect -3926 514574 -3306 514658
rect -3926 514338 -3894 514574
rect -3658 514338 -3574 514574
rect -3338 514338 -3306 514574
rect -3926 478894 -3306 514338
rect -3926 478658 -3894 478894
rect -3658 478658 -3574 478894
rect -3338 478658 -3306 478894
rect -3926 478574 -3306 478658
rect -3926 478338 -3894 478574
rect -3658 478338 -3574 478574
rect -3338 478338 -3306 478574
rect -3926 442894 -3306 478338
rect -3926 442658 -3894 442894
rect -3658 442658 -3574 442894
rect -3338 442658 -3306 442894
rect -3926 442574 -3306 442658
rect -3926 442338 -3894 442574
rect -3658 442338 -3574 442574
rect -3338 442338 -3306 442574
rect -3926 406894 -3306 442338
rect -3926 406658 -3894 406894
rect -3658 406658 -3574 406894
rect -3338 406658 -3306 406894
rect -3926 406574 -3306 406658
rect -3926 406338 -3894 406574
rect -3658 406338 -3574 406574
rect -3338 406338 -3306 406574
rect -3926 370894 -3306 406338
rect -3926 370658 -3894 370894
rect -3658 370658 -3574 370894
rect -3338 370658 -3306 370894
rect -3926 370574 -3306 370658
rect -3926 370338 -3894 370574
rect -3658 370338 -3574 370574
rect -3338 370338 -3306 370574
rect -3926 334894 -3306 370338
rect -3926 334658 -3894 334894
rect -3658 334658 -3574 334894
rect -3338 334658 -3306 334894
rect -3926 334574 -3306 334658
rect -3926 334338 -3894 334574
rect -3658 334338 -3574 334574
rect -3338 334338 -3306 334574
rect -3926 298894 -3306 334338
rect -3926 298658 -3894 298894
rect -3658 298658 -3574 298894
rect -3338 298658 -3306 298894
rect -3926 298574 -3306 298658
rect -3926 298338 -3894 298574
rect -3658 298338 -3574 298574
rect -3338 298338 -3306 298574
rect -3926 262894 -3306 298338
rect -3926 262658 -3894 262894
rect -3658 262658 -3574 262894
rect -3338 262658 -3306 262894
rect -3926 262574 -3306 262658
rect -3926 262338 -3894 262574
rect -3658 262338 -3574 262574
rect -3338 262338 -3306 262574
rect -3926 226894 -3306 262338
rect -3926 226658 -3894 226894
rect -3658 226658 -3574 226894
rect -3338 226658 -3306 226894
rect -3926 226574 -3306 226658
rect -3926 226338 -3894 226574
rect -3658 226338 -3574 226574
rect -3338 226338 -3306 226574
rect -3926 190894 -3306 226338
rect -3926 190658 -3894 190894
rect -3658 190658 -3574 190894
rect -3338 190658 -3306 190894
rect -3926 190574 -3306 190658
rect -3926 190338 -3894 190574
rect -3658 190338 -3574 190574
rect -3338 190338 -3306 190574
rect -3926 154894 -3306 190338
rect -3926 154658 -3894 154894
rect -3658 154658 -3574 154894
rect -3338 154658 -3306 154894
rect -3926 154574 -3306 154658
rect -3926 154338 -3894 154574
rect -3658 154338 -3574 154574
rect -3338 154338 -3306 154574
rect -3926 118894 -3306 154338
rect -3926 118658 -3894 118894
rect -3658 118658 -3574 118894
rect -3338 118658 -3306 118894
rect -3926 118574 -3306 118658
rect -3926 118338 -3894 118574
rect -3658 118338 -3574 118574
rect -3338 118338 -3306 118574
rect -3926 82894 -3306 118338
rect -3926 82658 -3894 82894
rect -3658 82658 -3574 82894
rect -3338 82658 -3306 82894
rect -3926 82574 -3306 82658
rect -3926 82338 -3894 82574
rect -3658 82338 -3574 82574
rect -3338 82338 -3306 82574
rect -3926 46894 -3306 82338
rect -3926 46658 -3894 46894
rect -3658 46658 -3574 46894
rect -3338 46658 -3306 46894
rect -3926 46574 -3306 46658
rect -3926 46338 -3894 46574
rect -3658 46338 -3574 46574
rect -3338 46338 -3306 46574
rect -3926 10894 -3306 46338
rect -3926 10658 -3894 10894
rect -3658 10658 -3574 10894
rect -3338 10658 -3306 10894
rect -3926 10574 -3306 10658
rect -3926 10338 -3894 10574
rect -3658 10338 -3574 10574
rect -3338 10338 -3306 10574
rect -3926 -2266 -3306 10338
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691174 -2346 705242
rect -2966 690938 -2934 691174
rect -2698 690938 -2614 691174
rect -2378 690938 -2346 691174
rect -2966 690854 -2346 690938
rect -2966 690618 -2934 690854
rect -2698 690618 -2614 690854
rect -2378 690618 -2346 690854
rect -2966 655174 -2346 690618
rect -2966 654938 -2934 655174
rect -2698 654938 -2614 655174
rect -2378 654938 -2346 655174
rect -2966 654854 -2346 654938
rect -2966 654618 -2934 654854
rect -2698 654618 -2614 654854
rect -2378 654618 -2346 654854
rect -2966 619174 -2346 654618
rect -2966 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 -2346 619174
rect -2966 618854 -2346 618938
rect -2966 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 -2346 618854
rect -2966 583174 -2346 618618
rect -2966 582938 -2934 583174
rect -2698 582938 -2614 583174
rect -2378 582938 -2346 583174
rect -2966 582854 -2346 582938
rect -2966 582618 -2934 582854
rect -2698 582618 -2614 582854
rect -2378 582618 -2346 582854
rect -2966 547174 -2346 582618
rect -2966 546938 -2934 547174
rect -2698 546938 -2614 547174
rect -2378 546938 -2346 547174
rect -2966 546854 -2346 546938
rect -2966 546618 -2934 546854
rect -2698 546618 -2614 546854
rect -2378 546618 -2346 546854
rect -2966 511174 -2346 546618
rect -2966 510938 -2934 511174
rect -2698 510938 -2614 511174
rect -2378 510938 -2346 511174
rect -2966 510854 -2346 510938
rect -2966 510618 -2934 510854
rect -2698 510618 -2614 510854
rect -2378 510618 -2346 510854
rect -2966 475174 -2346 510618
rect -2966 474938 -2934 475174
rect -2698 474938 -2614 475174
rect -2378 474938 -2346 475174
rect -2966 474854 -2346 474938
rect -2966 474618 -2934 474854
rect -2698 474618 -2614 474854
rect -2378 474618 -2346 474854
rect -2966 439174 -2346 474618
rect -2966 438938 -2934 439174
rect -2698 438938 -2614 439174
rect -2378 438938 -2346 439174
rect -2966 438854 -2346 438938
rect -2966 438618 -2934 438854
rect -2698 438618 -2614 438854
rect -2378 438618 -2346 438854
rect -2966 403174 -2346 438618
rect -2966 402938 -2934 403174
rect -2698 402938 -2614 403174
rect -2378 402938 -2346 403174
rect -2966 402854 -2346 402938
rect -2966 402618 -2934 402854
rect -2698 402618 -2614 402854
rect -2378 402618 -2346 402854
rect -2966 367174 -2346 402618
rect -2966 366938 -2934 367174
rect -2698 366938 -2614 367174
rect -2378 366938 -2346 367174
rect -2966 366854 -2346 366938
rect -2966 366618 -2934 366854
rect -2698 366618 -2614 366854
rect -2378 366618 -2346 366854
rect -2966 331174 -2346 366618
rect -2966 330938 -2934 331174
rect -2698 330938 -2614 331174
rect -2378 330938 -2346 331174
rect -2966 330854 -2346 330938
rect -2966 330618 -2934 330854
rect -2698 330618 -2614 330854
rect -2378 330618 -2346 330854
rect -2966 295174 -2346 330618
rect -2966 294938 -2934 295174
rect -2698 294938 -2614 295174
rect -2378 294938 -2346 295174
rect -2966 294854 -2346 294938
rect -2966 294618 -2934 294854
rect -2698 294618 -2614 294854
rect -2378 294618 -2346 294854
rect -2966 259174 -2346 294618
rect -2966 258938 -2934 259174
rect -2698 258938 -2614 259174
rect -2378 258938 -2346 259174
rect -2966 258854 -2346 258938
rect -2966 258618 -2934 258854
rect -2698 258618 -2614 258854
rect -2378 258618 -2346 258854
rect -2966 223174 -2346 258618
rect -2966 222938 -2934 223174
rect -2698 222938 -2614 223174
rect -2378 222938 -2346 223174
rect -2966 222854 -2346 222938
rect -2966 222618 -2934 222854
rect -2698 222618 -2614 222854
rect -2378 222618 -2346 222854
rect -2966 187174 -2346 222618
rect -2966 186938 -2934 187174
rect -2698 186938 -2614 187174
rect -2378 186938 -2346 187174
rect -2966 186854 -2346 186938
rect -2966 186618 -2934 186854
rect -2698 186618 -2614 186854
rect -2378 186618 -2346 186854
rect -2966 151174 -2346 186618
rect -2966 150938 -2934 151174
rect -2698 150938 -2614 151174
rect -2378 150938 -2346 151174
rect -2966 150854 -2346 150938
rect -2966 150618 -2934 150854
rect -2698 150618 -2614 150854
rect -2378 150618 -2346 150854
rect -2966 115174 -2346 150618
rect -2966 114938 -2934 115174
rect -2698 114938 -2614 115174
rect -2378 114938 -2346 115174
rect -2966 114854 -2346 114938
rect -2966 114618 -2934 114854
rect -2698 114618 -2614 114854
rect -2378 114618 -2346 114854
rect -2966 79174 -2346 114618
rect -2966 78938 -2934 79174
rect -2698 78938 -2614 79174
rect -2378 78938 -2346 79174
rect -2966 78854 -2346 78938
rect -2966 78618 -2934 78854
rect -2698 78618 -2614 78854
rect -2378 78618 -2346 78854
rect -2966 43174 -2346 78618
rect -2966 42938 -2934 43174
rect -2698 42938 -2614 43174
rect -2378 42938 -2346 43174
rect -2966 42854 -2346 42938
rect -2966 42618 -2934 42854
rect -2698 42618 -2614 42854
rect -2378 42618 -2346 42854
rect -2966 7174 -2346 42618
rect -2966 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 -2346 7174
rect -2966 6854 -2346 6938
rect -2966 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 -2346 6854
rect -2966 -1306 -2346 6618
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 9234 706758 9854 711590
rect 9234 706522 9266 706758
rect 9502 706522 9586 706758
rect 9822 706522 9854 706758
rect 9234 706438 9854 706522
rect 9234 706202 9266 706438
rect 9502 706202 9586 706438
rect 9822 706202 9854 706438
rect 9234 694894 9854 706202
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 692105 9854 694338
rect 12954 707718 13574 711590
rect 12954 707482 12986 707718
rect 13222 707482 13306 707718
rect 13542 707482 13574 707718
rect 12954 707398 13574 707482
rect 12954 707162 12986 707398
rect 13222 707162 13306 707398
rect 13542 707162 13574 707398
rect 12954 698614 13574 707162
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 692105 13574 698058
rect 45234 706758 45854 711590
rect 45234 706522 45266 706758
rect 45502 706522 45586 706758
rect 45822 706522 45854 706758
rect 45234 706438 45854 706522
rect 45234 706202 45266 706438
rect 45502 706202 45586 706438
rect 45822 706202 45854 706438
rect 45234 694894 45854 706202
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 692105 45854 694338
rect 48954 707718 49574 711590
rect 48954 707482 48986 707718
rect 49222 707482 49306 707718
rect 49542 707482 49574 707718
rect 48954 707398 49574 707482
rect 48954 707162 48986 707398
rect 49222 707162 49306 707398
rect 49542 707162 49574 707398
rect 48954 698614 49574 707162
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 692105 49574 698058
rect 81234 706758 81854 711590
rect 81234 706522 81266 706758
rect 81502 706522 81586 706758
rect 81822 706522 81854 706758
rect 81234 706438 81854 706522
rect 81234 706202 81266 706438
rect 81502 706202 81586 706438
rect 81822 706202 81854 706438
rect 81234 694894 81854 706202
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 692105 81854 694338
rect 84954 707718 85574 711590
rect 84954 707482 84986 707718
rect 85222 707482 85306 707718
rect 85542 707482 85574 707718
rect 84954 707398 85574 707482
rect 84954 707162 84986 707398
rect 85222 707162 85306 707398
rect 85542 707162 85574 707398
rect 84954 698614 85574 707162
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 692105 85574 698058
rect 117234 706758 117854 711590
rect 117234 706522 117266 706758
rect 117502 706522 117586 706758
rect 117822 706522 117854 706758
rect 117234 706438 117854 706522
rect 117234 706202 117266 706438
rect 117502 706202 117586 706438
rect 117822 706202 117854 706438
rect 117234 694894 117854 706202
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 692460 117854 694338
rect 120954 707718 121574 711590
rect 120954 707482 120986 707718
rect 121222 707482 121306 707718
rect 121542 707482 121574 707718
rect 120954 707398 121574 707482
rect 120954 707162 120986 707398
rect 121222 707162 121306 707398
rect 121542 707162 121574 707398
rect 120954 698614 121574 707162
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 692105 121574 698058
rect 153234 706758 153854 711590
rect 153234 706522 153266 706758
rect 153502 706522 153586 706758
rect 153822 706522 153854 706758
rect 153234 706438 153854 706522
rect 153234 706202 153266 706438
rect 153502 706202 153586 706438
rect 153822 706202 153854 706438
rect 153234 694894 153854 706202
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 692105 153854 694338
rect 156954 707718 157574 711590
rect 156954 707482 156986 707718
rect 157222 707482 157306 707718
rect 157542 707482 157574 707718
rect 156954 707398 157574 707482
rect 156954 707162 156986 707398
rect 157222 707162 157306 707398
rect 157542 707162 157574 707398
rect 156954 698614 157574 707162
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 692105 157574 698058
rect 189234 706758 189854 711590
rect 189234 706522 189266 706758
rect 189502 706522 189586 706758
rect 189822 706522 189854 706758
rect 189234 706438 189854 706522
rect 189234 706202 189266 706438
rect 189502 706202 189586 706438
rect 189822 706202 189854 706438
rect 189234 694894 189854 706202
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 692105 189854 694338
rect 192954 707718 193574 711590
rect 192954 707482 192986 707718
rect 193222 707482 193306 707718
rect 193542 707482 193574 707718
rect 192954 707398 193574 707482
rect 192954 707162 192986 707398
rect 193222 707162 193306 707398
rect 193542 707162 193574 707398
rect 192954 698614 193574 707162
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 692105 193574 698058
rect 225234 706758 225854 711590
rect 225234 706522 225266 706758
rect 225502 706522 225586 706758
rect 225822 706522 225854 706758
rect 225234 706438 225854 706522
rect 225234 706202 225266 706438
rect 225502 706202 225586 706438
rect 225822 706202 225854 706438
rect 225234 694894 225854 706202
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 692460 225854 694338
rect 228954 707718 229574 711590
rect 228954 707482 228986 707718
rect 229222 707482 229306 707718
rect 229542 707482 229574 707718
rect 228954 707398 229574 707482
rect 228954 707162 228986 707398
rect 229222 707162 229306 707398
rect 229542 707162 229574 707398
rect 228954 698614 229574 707162
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 692105 229574 698058
rect 261234 706758 261854 711590
rect 261234 706522 261266 706758
rect 261502 706522 261586 706758
rect 261822 706522 261854 706758
rect 261234 706438 261854 706522
rect 261234 706202 261266 706438
rect 261502 706202 261586 706438
rect 261822 706202 261854 706438
rect 261234 694894 261854 706202
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 692105 261854 694338
rect 264954 707718 265574 711590
rect 264954 707482 264986 707718
rect 265222 707482 265306 707718
rect 265542 707482 265574 707718
rect 264954 707398 265574 707482
rect 264954 707162 264986 707398
rect 265222 707162 265306 707398
rect 265542 707162 265574 707398
rect 264954 698614 265574 707162
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 692105 265574 698058
rect 297234 706758 297854 711590
rect 297234 706522 297266 706758
rect 297502 706522 297586 706758
rect 297822 706522 297854 706758
rect 297234 706438 297854 706522
rect 297234 706202 297266 706438
rect 297502 706202 297586 706438
rect 297822 706202 297854 706438
rect 297234 694894 297854 706202
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 692105 297854 694338
rect 300954 707718 301574 711590
rect 300954 707482 300986 707718
rect 301222 707482 301306 707718
rect 301542 707482 301574 707718
rect 300954 707398 301574 707482
rect 300954 707162 300986 707398
rect 301222 707162 301306 707398
rect 301542 707162 301574 707398
rect 300954 698614 301574 707162
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 692105 301574 698058
rect 333234 706758 333854 711590
rect 333234 706522 333266 706758
rect 333502 706522 333586 706758
rect 333822 706522 333854 706758
rect 333234 706438 333854 706522
rect 333234 706202 333266 706438
rect 333502 706202 333586 706438
rect 333822 706202 333854 706438
rect 333234 694894 333854 706202
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 692105 333854 694338
rect 336954 707718 337574 711590
rect 336954 707482 336986 707718
rect 337222 707482 337306 707718
rect 337542 707482 337574 707718
rect 336954 707398 337574 707482
rect 336954 707162 336986 707398
rect 337222 707162 337306 707398
rect 337542 707162 337574 707398
rect 336954 698614 337574 707162
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 692105 337574 698058
rect 369234 706758 369854 711590
rect 369234 706522 369266 706758
rect 369502 706522 369586 706758
rect 369822 706522 369854 706758
rect 369234 706438 369854 706522
rect 369234 706202 369266 706438
rect 369502 706202 369586 706438
rect 369822 706202 369854 706438
rect 369234 694894 369854 706202
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 692105 369854 694338
rect 372954 707718 373574 711590
rect 372954 707482 372986 707718
rect 373222 707482 373306 707718
rect 373542 707482 373574 707718
rect 372954 707398 373574 707482
rect 372954 707162 372986 707398
rect 373222 707162 373306 707398
rect 373542 707162 373574 707398
rect 372954 698614 373574 707162
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 692105 373574 698058
rect 405234 706758 405854 711590
rect 405234 706522 405266 706758
rect 405502 706522 405586 706758
rect 405822 706522 405854 706758
rect 405234 706438 405854 706522
rect 405234 706202 405266 706438
rect 405502 706202 405586 706438
rect 405822 706202 405854 706438
rect 405234 694894 405854 706202
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 692105 405854 694338
rect 408954 707718 409574 711590
rect 408954 707482 408986 707718
rect 409222 707482 409306 707718
rect 409542 707482 409574 707718
rect 408954 707398 409574 707482
rect 408954 707162 408986 707398
rect 409222 707162 409306 707398
rect 409542 707162 409574 707398
rect 408954 698614 409574 707162
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 692460 409574 698058
rect 441234 706758 441854 711590
rect 441234 706522 441266 706758
rect 441502 706522 441586 706758
rect 441822 706522 441854 706758
rect 441234 706438 441854 706522
rect 441234 706202 441266 706438
rect 441502 706202 441586 706438
rect 441822 706202 441854 706438
rect 441234 694894 441854 706202
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 692105 441854 694338
rect 444954 707718 445574 711590
rect 444954 707482 444986 707718
rect 445222 707482 445306 707718
rect 445542 707482 445574 707718
rect 444954 707398 445574 707482
rect 444954 707162 444986 707398
rect 445222 707162 445306 707398
rect 445542 707162 445574 707398
rect 444954 698614 445574 707162
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 692105 445574 698058
rect 477234 706758 477854 711590
rect 477234 706522 477266 706758
rect 477502 706522 477586 706758
rect 477822 706522 477854 706758
rect 477234 706438 477854 706522
rect 477234 706202 477266 706438
rect 477502 706202 477586 706438
rect 477822 706202 477854 706438
rect 477234 694894 477854 706202
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 692105 477854 694338
rect 480954 707718 481574 711590
rect 480954 707482 480986 707718
rect 481222 707482 481306 707718
rect 481542 707482 481574 707718
rect 480954 707398 481574 707482
rect 480954 707162 480986 707398
rect 481222 707162 481306 707398
rect 481542 707162 481574 707398
rect 480954 698614 481574 707162
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 692105 481574 698058
rect 513234 706758 513854 711590
rect 513234 706522 513266 706758
rect 513502 706522 513586 706758
rect 513822 706522 513854 706758
rect 513234 706438 513854 706522
rect 513234 706202 513266 706438
rect 513502 706202 513586 706438
rect 513822 706202 513854 706438
rect 513234 694894 513854 706202
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 692105 513854 694338
rect 516954 707718 517574 711590
rect 516954 707482 516986 707718
rect 517222 707482 517306 707718
rect 517542 707482 517574 707718
rect 516954 707398 517574 707482
rect 516954 707162 516986 707398
rect 517222 707162 517306 707398
rect 517542 707162 517574 707398
rect 516954 698614 517574 707162
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 692460 517574 698058
rect 549234 706758 549854 711590
rect 549234 706522 549266 706758
rect 549502 706522 549586 706758
rect 549822 706522 549854 706758
rect 549234 706438 549854 706522
rect 549234 706202 549266 706438
rect 549502 706202 549586 706438
rect 549822 706202 549854 706438
rect 549234 694894 549854 706202
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 692105 549854 694338
rect 552954 707718 553574 711590
rect 552954 707482 552986 707718
rect 553222 707482 553306 707718
rect 553542 707482 553574 707718
rect 552954 707398 553574 707482
rect 552954 707162 552986 707398
rect 553222 707162 553306 707398
rect 553542 707162 553574 707398
rect 552954 698614 553574 707162
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 692105 553574 698058
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 10208 687454 10528 687486
rect 10208 687218 10250 687454
rect 10486 687218 10528 687454
rect 10208 687134 10528 687218
rect 10208 686898 10250 687134
rect 10486 686898 10528 687134
rect 10208 686866 10528 686898
rect 40928 687454 41248 687486
rect 40928 687218 40970 687454
rect 41206 687218 41248 687454
rect 40928 687134 41248 687218
rect 40928 686898 40970 687134
rect 41206 686898 41248 687134
rect 40928 686866 41248 686898
rect 71648 687454 71968 687486
rect 71648 687218 71690 687454
rect 71926 687218 71968 687454
rect 71648 687134 71968 687218
rect 71648 686898 71690 687134
rect 71926 686898 71968 687134
rect 71648 686866 71968 686898
rect 102368 687454 102688 687486
rect 102368 687218 102410 687454
rect 102646 687218 102688 687454
rect 102368 687134 102688 687218
rect 102368 686898 102410 687134
rect 102646 686898 102688 687134
rect 102368 686866 102688 686898
rect 133088 687454 133408 687486
rect 133088 687218 133130 687454
rect 133366 687218 133408 687454
rect 133088 687134 133408 687218
rect 133088 686898 133130 687134
rect 133366 686898 133408 687134
rect 133088 686866 133408 686898
rect 163808 687454 164128 687486
rect 163808 687218 163850 687454
rect 164086 687218 164128 687454
rect 163808 687134 164128 687218
rect 163808 686898 163850 687134
rect 164086 686898 164128 687134
rect 163808 686866 164128 686898
rect 194528 687454 194848 687486
rect 194528 687218 194570 687454
rect 194806 687218 194848 687454
rect 194528 687134 194848 687218
rect 194528 686898 194570 687134
rect 194806 686898 194848 687134
rect 194528 686866 194848 686898
rect 225248 687454 225568 687486
rect 225248 687218 225290 687454
rect 225526 687218 225568 687454
rect 225248 687134 225568 687218
rect 225248 686898 225290 687134
rect 225526 686898 225568 687134
rect 225248 686866 225568 686898
rect 255968 687454 256288 687486
rect 255968 687218 256010 687454
rect 256246 687218 256288 687454
rect 255968 687134 256288 687218
rect 255968 686898 256010 687134
rect 256246 686898 256288 687134
rect 255968 686866 256288 686898
rect 286688 687454 287008 687486
rect 286688 687218 286730 687454
rect 286966 687218 287008 687454
rect 286688 687134 287008 687218
rect 286688 686898 286730 687134
rect 286966 686898 287008 687134
rect 286688 686866 287008 686898
rect 317408 687454 317728 687486
rect 317408 687218 317450 687454
rect 317686 687218 317728 687454
rect 317408 687134 317728 687218
rect 317408 686898 317450 687134
rect 317686 686898 317728 687134
rect 317408 686866 317728 686898
rect 348128 687454 348448 687486
rect 348128 687218 348170 687454
rect 348406 687218 348448 687454
rect 348128 687134 348448 687218
rect 348128 686898 348170 687134
rect 348406 686898 348448 687134
rect 348128 686866 348448 686898
rect 378848 687454 379168 687486
rect 378848 687218 378890 687454
rect 379126 687218 379168 687454
rect 378848 687134 379168 687218
rect 378848 686898 378890 687134
rect 379126 686898 379168 687134
rect 378848 686866 379168 686898
rect 409568 687454 409888 687486
rect 409568 687218 409610 687454
rect 409846 687218 409888 687454
rect 409568 687134 409888 687218
rect 409568 686898 409610 687134
rect 409846 686898 409888 687134
rect 409568 686866 409888 686898
rect 440288 687454 440608 687486
rect 440288 687218 440330 687454
rect 440566 687218 440608 687454
rect 440288 687134 440608 687218
rect 440288 686898 440330 687134
rect 440566 686898 440608 687134
rect 440288 686866 440608 686898
rect 471008 687454 471328 687486
rect 471008 687218 471050 687454
rect 471286 687218 471328 687454
rect 471008 687134 471328 687218
rect 471008 686898 471050 687134
rect 471286 686898 471328 687134
rect 471008 686866 471328 686898
rect 501728 687454 502048 687486
rect 501728 687218 501770 687454
rect 502006 687218 502048 687454
rect 501728 687134 502048 687218
rect 501728 686898 501770 687134
rect 502006 686898 502048 687134
rect 501728 686866 502048 686898
rect 532448 687454 532768 687486
rect 532448 687218 532490 687454
rect 532726 687218 532768 687454
rect 532448 687134 532768 687218
rect 532448 686898 532490 687134
rect 532726 686898 532768 687134
rect 532448 686866 532768 686898
rect 563168 687454 563488 687486
rect 563168 687218 563210 687454
rect 563446 687218 563488 687454
rect 563168 687134 563488 687218
rect 563168 686898 563210 687134
rect 563446 686898 563488 687134
rect 563168 686866 563488 686898
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 25568 655174 25888 655206
rect 25568 654938 25610 655174
rect 25846 654938 25888 655174
rect 25568 654854 25888 654938
rect 25568 654618 25610 654854
rect 25846 654618 25888 654854
rect 25568 654586 25888 654618
rect 56288 655174 56608 655206
rect 56288 654938 56330 655174
rect 56566 654938 56608 655174
rect 56288 654854 56608 654938
rect 56288 654618 56330 654854
rect 56566 654618 56608 654854
rect 56288 654586 56608 654618
rect 87008 655174 87328 655206
rect 87008 654938 87050 655174
rect 87286 654938 87328 655174
rect 87008 654854 87328 654938
rect 87008 654618 87050 654854
rect 87286 654618 87328 654854
rect 87008 654586 87328 654618
rect 117728 655174 118048 655206
rect 117728 654938 117770 655174
rect 118006 654938 118048 655174
rect 117728 654854 118048 654938
rect 117728 654618 117770 654854
rect 118006 654618 118048 654854
rect 117728 654586 118048 654618
rect 148448 655174 148768 655206
rect 148448 654938 148490 655174
rect 148726 654938 148768 655174
rect 148448 654854 148768 654938
rect 148448 654618 148490 654854
rect 148726 654618 148768 654854
rect 148448 654586 148768 654618
rect 179168 655174 179488 655206
rect 179168 654938 179210 655174
rect 179446 654938 179488 655174
rect 179168 654854 179488 654938
rect 179168 654618 179210 654854
rect 179446 654618 179488 654854
rect 179168 654586 179488 654618
rect 209888 655174 210208 655206
rect 209888 654938 209930 655174
rect 210166 654938 210208 655174
rect 209888 654854 210208 654938
rect 209888 654618 209930 654854
rect 210166 654618 210208 654854
rect 209888 654586 210208 654618
rect 240608 655174 240928 655206
rect 240608 654938 240650 655174
rect 240886 654938 240928 655174
rect 240608 654854 240928 654938
rect 240608 654618 240650 654854
rect 240886 654618 240928 654854
rect 240608 654586 240928 654618
rect 271328 655174 271648 655206
rect 271328 654938 271370 655174
rect 271606 654938 271648 655174
rect 271328 654854 271648 654938
rect 271328 654618 271370 654854
rect 271606 654618 271648 654854
rect 271328 654586 271648 654618
rect 302048 655174 302368 655206
rect 302048 654938 302090 655174
rect 302326 654938 302368 655174
rect 302048 654854 302368 654938
rect 302048 654618 302090 654854
rect 302326 654618 302368 654854
rect 302048 654586 302368 654618
rect 332768 655174 333088 655206
rect 332768 654938 332810 655174
rect 333046 654938 333088 655174
rect 332768 654854 333088 654938
rect 332768 654618 332810 654854
rect 333046 654618 333088 654854
rect 332768 654586 333088 654618
rect 363488 655174 363808 655206
rect 363488 654938 363530 655174
rect 363766 654938 363808 655174
rect 363488 654854 363808 654938
rect 363488 654618 363530 654854
rect 363766 654618 363808 654854
rect 363488 654586 363808 654618
rect 394208 655174 394528 655206
rect 394208 654938 394250 655174
rect 394486 654938 394528 655174
rect 394208 654854 394528 654938
rect 394208 654618 394250 654854
rect 394486 654618 394528 654854
rect 394208 654586 394528 654618
rect 424928 655174 425248 655206
rect 424928 654938 424970 655174
rect 425206 654938 425248 655174
rect 424928 654854 425248 654938
rect 424928 654618 424970 654854
rect 425206 654618 425248 654854
rect 424928 654586 425248 654618
rect 455648 655174 455968 655206
rect 455648 654938 455690 655174
rect 455926 654938 455968 655174
rect 455648 654854 455968 654938
rect 455648 654618 455690 654854
rect 455926 654618 455968 654854
rect 455648 654586 455968 654618
rect 486368 655174 486688 655206
rect 486368 654938 486410 655174
rect 486646 654938 486688 655174
rect 486368 654854 486688 654938
rect 486368 654618 486410 654854
rect 486646 654618 486688 654854
rect 486368 654586 486688 654618
rect 517088 655174 517408 655206
rect 517088 654938 517130 655174
rect 517366 654938 517408 655174
rect 517088 654854 517408 654938
rect 517088 654618 517130 654854
rect 517366 654618 517408 654854
rect 517088 654586 517408 654618
rect 547808 655174 548128 655206
rect 547808 654938 547850 655174
rect 548086 654938 548128 655174
rect 547808 654854 548128 654938
rect 547808 654618 547850 654854
rect 548086 654618 548128 654854
rect 547808 654586 548128 654618
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 10208 651454 10528 651486
rect 10208 651218 10250 651454
rect 10486 651218 10528 651454
rect 10208 651134 10528 651218
rect 10208 650898 10250 651134
rect 10486 650898 10528 651134
rect 10208 650866 10528 650898
rect 40928 651454 41248 651486
rect 40928 651218 40970 651454
rect 41206 651218 41248 651454
rect 40928 651134 41248 651218
rect 40928 650898 40970 651134
rect 41206 650898 41248 651134
rect 40928 650866 41248 650898
rect 71648 651454 71968 651486
rect 71648 651218 71690 651454
rect 71926 651218 71968 651454
rect 71648 651134 71968 651218
rect 71648 650898 71690 651134
rect 71926 650898 71968 651134
rect 71648 650866 71968 650898
rect 102368 651454 102688 651486
rect 102368 651218 102410 651454
rect 102646 651218 102688 651454
rect 102368 651134 102688 651218
rect 102368 650898 102410 651134
rect 102646 650898 102688 651134
rect 102368 650866 102688 650898
rect 133088 651454 133408 651486
rect 133088 651218 133130 651454
rect 133366 651218 133408 651454
rect 133088 651134 133408 651218
rect 133088 650898 133130 651134
rect 133366 650898 133408 651134
rect 133088 650866 133408 650898
rect 163808 651454 164128 651486
rect 163808 651218 163850 651454
rect 164086 651218 164128 651454
rect 163808 651134 164128 651218
rect 163808 650898 163850 651134
rect 164086 650898 164128 651134
rect 163808 650866 164128 650898
rect 194528 651454 194848 651486
rect 194528 651218 194570 651454
rect 194806 651218 194848 651454
rect 194528 651134 194848 651218
rect 194528 650898 194570 651134
rect 194806 650898 194848 651134
rect 194528 650866 194848 650898
rect 225248 651454 225568 651486
rect 225248 651218 225290 651454
rect 225526 651218 225568 651454
rect 225248 651134 225568 651218
rect 225248 650898 225290 651134
rect 225526 650898 225568 651134
rect 225248 650866 225568 650898
rect 255968 651454 256288 651486
rect 255968 651218 256010 651454
rect 256246 651218 256288 651454
rect 255968 651134 256288 651218
rect 255968 650898 256010 651134
rect 256246 650898 256288 651134
rect 255968 650866 256288 650898
rect 286688 651454 287008 651486
rect 286688 651218 286730 651454
rect 286966 651218 287008 651454
rect 286688 651134 287008 651218
rect 286688 650898 286730 651134
rect 286966 650898 287008 651134
rect 286688 650866 287008 650898
rect 317408 651454 317728 651486
rect 317408 651218 317450 651454
rect 317686 651218 317728 651454
rect 317408 651134 317728 651218
rect 317408 650898 317450 651134
rect 317686 650898 317728 651134
rect 317408 650866 317728 650898
rect 348128 651454 348448 651486
rect 348128 651218 348170 651454
rect 348406 651218 348448 651454
rect 348128 651134 348448 651218
rect 348128 650898 348170 651134
rect 348406 650898 348448 651134
rect 348128 650866 348448 650898
rect 378848 651454 379168 651486
rect 378848 651218 378890 651454
rect 379126 651218 379168 651454
rect 378848 651134 379168 651218
rect 378848 650898 378890 651134
rect 379126 650898 379168 651134
rect 378848 650866 379168 650898
rect 409568 651454 409888 651486
rect 409568 651218 409610 651454
rect 409846 651218 409888 651454
rect 409568 651134 409888 651218
rect 409568 650898 409610 651134
rect 409846 650898 409888 651134
rect 409568 650866 409888 650898
rect 440288 651454 440608 651486
rect 440288 651218 440330 651454
rect 440566 651218 440608 651454
rect 440288 651134 440608 651218
rect 440288 650898 440330 651134
rect 440566 650898 440608 651134
rect 440288 650866 440608 650898
rect 471008 651454 471328 651486
rect 471008 651218 471050 651454
rect 471286 651218 471328 651454
rect 471008 651134 471328 651218
rect 471008 650898 471050 651134
rect 471286 650898 471328 651134
rect 471008 650866 471328 650898
rect 501728 651454 502048 651486
rect 501728 651218 501770 651454
rect 502006 651218 502048 651454
rect 501728 651134 502048 651218
rect 501728 650898 501770 651134
rect 502006 650898 502048 651134
rect 501728 650866 502048 650898
rect 532448 651454 532768 651486
rect 532448 651218 532490 651454
rect 532726 651218 532768 651454
rect 532448 651134 532768 651218
rect 532448 650898 532490 651134
rect 532726 650898 532768 651134
rect 532448 650866 532768 650898
rect 563168 651454 563488 651486
rect 563168 651218 563210 651454
rect 563446 651218 563488 651454
rect 563168 651134 563488 651218
rect 563168 650898 563210 651134
rect 563446 650898 563488 651134
rect 563168 650866 563488 650898
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 25568 619174 25888 619206
rect 25568 618938 25610 619174
rect 25846 618938 25888 619174
rect 25568 618854 25888 618938
rect 25568 618618 25610 618854
rect 25846 618618 25888 618854
rect 25568 618586 25888 618618
rect 56288 619174 56608 619206
rect 56288 618938 56330 619174
rect 56566 618938 56608 619174
rect 56288 618854 56608 618938
rect 56288 618618 56330 618854
rect 56566 618618 56608 618854
rect 56288 618586 56608 618618
rect 87008 619174 87328 619206
rect 87008 618938 87050 619174
rect 87286 618938 87328 619174
rect 87008 618854 87328 618938
rect 87008 618618 87050 618854
rect 87286 618618 87328 618854
rect 87008 618586 87328 618618
rect 117728 619174 118048 619206
rect 117728 618938 117770 619174
rect 118006 618938 118048 619174
rect 117728 618854 118048 618938
rect 117728 618618 117770 618854
rect 118006 618618 118048 618854
rect 117728 618586 118048 618618
rect 148448 619174 148768 619206
rect 148448 618938 148490 619174
rect 148726 618938 148768 619174
rect 148448 618854 148768 618938
rect 148448 618618 148490 618854
rect 148726 618618 148768 618854
rect 148448 618586 148768 618618
rect 179168 619174 179488 619206
rect 179168 618938 179210 619174
rect 179446 618938 179488 619174
rect 179168 618854 179488 618938
rect 179168 618618 179210 618854
rect 179446 618618 179488 618854
rect 179168 618586 179488 618618
rect 209888 619174 210208 619206
rect 209888 618938 209930 619174
rect 210166 618938 210208 619174
rect 209888 618854 210208 618938
rect 209888 618618 209930 618854
rect 210166 618618 210208 618854
rect 209888 618586 210208 618618
rect 240608 619174 240928 619206
rect 240608 618938 240650 619174
rect 240886 618938 240928 619174
rect 240608 618854 240928 618938
rect 240608 618618 240650 618854
rect 240886 618618 240928 618854
rect 240608 618586 240928 618618
rect 271328 619174 271648 619206
rect 271328 618938 271370 619174
rect 271606 618938 271648 619174
rect 271328 618854 271648 618938
rect 271328 618618 271370 618854
rect 271606 618618 271648 618854
rect 271328 618586 271648 618618
rect 302048 619174 302368 619206
rect 302048 618938 302090 619174
rect 302326 618938 302368 619174
rect 302048 618854 302368 618938
rect 302048 618618 302090 618854
rect 302326 618618 302368 618854
rect 302048 618586 302368 618618
rect 332768 619174 333088 619206
rect 332768 618938 332810 619174
rect 333046 618938 333088 619174
rect 332768 618854 333088 618938
rect 332768 618618 332810 618854
rect 333046 618618 333088 618854
rect 332768 618586 333088 618618
rect 363488 619174 363808 619206
rect 363488 618938 363530 619174
rect 363766 618938 363808 619174
rect 363488 618854 363808 618938
rect 363488 618618 363530 618854
rect 363766 618618 363808 618854
rect 363488 618586 363808 618618
rect 394208 619174 394528 619206
rect 394208 618938 394250 619174
rect 394486 618938 394528 619174
rect 394208 618854 394528 618938
rect 394208 618618 394250 618854
rect 394486 618618 394528 618854
rect 394208 618586 394528 618618
rect 424928 619174 425248 619206
rect 424928 618938 424970 619174
rect 425206 618938 425248 619174
rect 424928 618854 425248 618938
rect 424928 618618 424970 618854
rect 425206 618618 425248 618854
rect 424928 618586 425248 618618
rect 455648 619174 455968 619206
rect 455648 618938 455690 619174
rect 455926 618938 455968 619174
rect 455648 618854 455968 618938
rect 455648 618618 455690 618854
rect 455926 618618 455968 618854
rect 455648 618586 455968 618618
rect 486368 619174 486688 619206
rect 486368 618938 486410 619174
rect 486646 618938 486688 619174
rect 486368 618854 486688 618938
rect 486368 618618 486410 618854
rect 486646 618618 486688 618854
rect 486368 618586 486688 618618
rect 517088 619174 517408 619206
rect 517088 618938 517130 619174
rect 517366 618938 517408 619174
rect 517088 618854 517408 618938
rect 517088 618618 517130 618854
rect 517366 618618 517408 618854
rect 517088 618586 517408 618618
rect 547808 619174 548128 619206
rect 547808 618938 547850 619174
rect 548086 618938 548128 619174
rect 547808 618854 548128 618938
rect 547808 618618 547850 618854
rect 548086 618618 548128 618854
rect 547808 618586 548128 618618
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 10208 615454 10528 615486
rect 10208 615218 10250 615454
rect 10486 615218 10528 615454
rect 10208 615134 10528 615218
rect 10208 614898 10250 615134
rect 10486 614898 10528 615134
rect 10208 614866 10528 614898
rect 40928 615454 41248 615486
rect 40928 615218 40970 615454
rect 41206 615218 41248 615454
rect 40928 615134 41248 615218
rect 40928 614898 40970 615134
rect 41206 614898 41248 615134
rect 40928 614866 41248 614898
rect 71648 615454 71968 615486
rect 71648 615218 71690 615454
rect 71926 615218 71968 615454
rect 71648 615134 71968 615218
rect 71648 614898 71690 615134
rect 71926 614898 71968 615134
rect 71648 614866 71968 614898
rect 102368 615454 102688 615486
rect 102368 615218 102410 615454
rect 102646 615218 102688 615454
rect 102368 615134 102688 615218
rect 102368 614898 102410 615134
rect 102646 614898 102688 615134
rect 102368 614866 102688 614898
rect 133088 615454 133408 615486
rect 133088 615218 133130 615454
rect 133366 615218 133408 615454
rect 133088 615134 133408 615218
rect 133088 614898 133130 615134
rect 133366 614898 133408 615134
rect 133088 614866 133408 614898
rect 163808 615454 164128 615486
rect 163808 615218 163850 615454
rect 164086 615218 164128 615454
rect 163808 615134 164128 615218
rect 163808 614898 163850 615134
rect 164086 614898 164128 615134
rect 163808 614866 164128 614898
rect 194528 615454 194848 615486
rect 194528 615218 194570 615454
rect 194806 615218 194848 615454
rect 194528 615134 194848 615218
rect 194528 614898 194570 615134
rect 194806 614898 194848 615134
rect 194528 614866 194848 614898
rect 225248 615454 225568 615486
rect 225248 615218 225290 615454
rect 225526 615218 225568 615454
rect 225248 615134 225568 615218
rect 225248 614898 225290 615134
rect 225526 614898 225568 615134
rect 225248 614866 225568 614898
rect 255968 615454 256288 615486
rect 255968 615218 256010 615454
rect 256246 615218 256288 615454
rect 255968 615134 256288 615218
rect 255968 614898 256010 615134
rect 256246 614898 256288 615134
rect 255968 614866 256288 614898
rect 286688 615454 287008 615486
rect 286688 615218 286730 615454
rect 286966 615218 287008 615454
rect 286688 615134 287008 615218
rect 286688 614898 286730 615134
rect 286966 614898 287008 615134
rect 286688 614866 287008 614898
rect 317408 615454 317728 615486
rect 317408 615218 317450 615454
rect 317686 615218 317728 615454
rect 317408 615134 317728 615218
rect 317408 614898 317450 615134
rect 317686 614898 317728 615134
rect 317408 614866 317728 614898
rect 348128 615454 348448 615486
rect 348128 615218 348170 615454
rect 348406 615218 348448 615454
rect 348128 615134 348448 615218
rect 348128 614898 348170 615134
rect 348406 614898 348448 615134
rect 348128 614866 348448 614898
rect 378848 615454 379168 615486
rect 378848 615218 378890 615454
rect 379126 615218 379168 615454
rect 378848 615134 379168 615218
rect 378848 614898 378890 615134
rect 379126 614898 379168 615134
rect 378848 614866 379168 614898
rect 409568 615454 409888 615486
rect 409568 615218 409610 615454
rect 409846 615218 409888 615454
rect 409568 615134 409888 615218
rect 409568 614898 409610 615134
rect 409846 614898 409888 615134
rect 409568 614866 409888 614898
rect 440288 615454 440608 615486
rect 440288 615218 440330 615454
rect 440566 615218 440608 615454
rect 440288 615134 440608 615218
rect 440288 614898 440330 615134
rect 440566 614898 440608 615134
rect 440288 614866 440608 614898
rect 471008 615454 471328 615486
rect 471008 615218 471050 615454
rect 471286 615218 471328 615454
rect 471008 615134 471328 615218
rect 471008 614898 471050 615134
rect 471286 614898 471328 615134
rect 471008 614866 471328 614898
rect 501728 615454 502048 615486
rect 501728 615218 501770 615454
rect 502006 615218 502048 615454
rect 501728 615134 502048 615218
rect 501728 614898 501770 615134
rect 502006 614898 502048 615134
rect 501728 614866 502048 614898
rect 532448 615454 532768 615486
rect 532448 615218 532490 615454
rect 532726 615218 532768 615454
rect 532448 615134 532768 615218
rect 532448 614898 532490 615134
rect 532726 614898 532768 615134
rect 532448 614866 532768 614898
rect 563168 615454 563488 615486
rect 563168 615218 563210 615454
rect 563446 615218 563488 615454
rect 563168 615134 563488 615218
rect 563168 614898 563210 615134
rect 563446 614898 563488 615134
rect 563168 614866 563488 614898
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 25568 583174 25888 583206
rect 25568 582938 25610 583174
rect 25846 582938 25888 583174
rect 25568 582854 25888 582938
rect 25568 582618 25610 582854
rect 25846 582618 25888 582854
rect 25568 582586 25888 582618
rect 56288 583174 56608 583206
rect 56288 582938 56330 583174
rect 56566 582938 56608 583174
rect 56288 582854 56608 582938
rect 56288 582618 56330 582854
rect 56566 582618 56608 582854
rect 56288 582586 56608 582618
rect 87008 583174 87328 583206
rect 87008 582938 87050 583174
rect 87286 582938 87328 583174
rect 87008 582854 87328 582938
rect 87008 582618 87050 582854
rect 87286 582618 87328 582854
rect 87008 582586 87328 582618
rect 117728 583174 118048 583206
rect 117728 582938 117770 583174
rect 118006 582938 118048 583174
rect 117728 582854 118048 582938
rect 117728 582618 117770 582854
rect 118006 582618 118048 582854
rect 117728 582586 118048 582618
rect 148448 583174 148768 583206
rect 148448 582938 148490 583174
rect 148726 582938 148768 583174
rect 148448 582854 148768 582938
rect 148448 582618 148490 582854
rect 148726 582618 148768 582854
rect 148448 582586 148768 582618
rect 179168 583174 179488 583206
rect 179168 582938 179210 583174
rect 179446 582938 179488 583174
rect 179168 582854 179488 582938
rect 179168 582618 179210 582854
rect 179446 582618 179488 582854
rect 179168 582586 179488 582618
rect 209888 583174 210208 583206
rect 209888 582938 209930 583174
rect 210166 582938 210208 583174
rect 209888 582854 210208 582938
rect 209888 582618 209930 582854
rect 210166 582618 210208 582854
rect 209888 582586 210208 582618
rect 240608 583174 240928 583206
rect 240608 582938 240650 583174
rect 240886 582938 240928 583174
rect 240608 582854 240928 582938
rect 240608 582618 240650 582854
rect 240886 582618 240928 582854
rect 240608 582586 240928 582618
rect 271328 583174 271648 583206
rect 271328 582938 271370 583174
rect 271606 582938 271648 583174
rect 271328 582854 271648 582938
rect 271328 582618 271370 582854
rect 271606 582618 271648 582854
rect 271328 582586 271648 582618
rect 302048 583174 302368 583206
rect 302048 582938 302090 583174
rect 302326 582938 302368 583174
rect 302048 582854 302368 582938
rect 302048 582618 302090 582854
rect 302326 582618 302368 582854
rect 302048 582586 302368 582618
rect 332768 583174 333088 583206
rect 332768 582938 332810 583174
rect 333046 582938 333088 583174
rect 332768 582854 333088 582938
rect 332768 582618 332810 582854
rect 333046 582618 333088 582854
rect 332768 582586 333088 582618
rect 363488 583174 363808 583206
rect 363488 582938 363530 583174
rect 363766 582938 363808 583174
rect 363488 582854 363808 582938
rect 363488 582618 363530 582854
rect 363766 582618 363808 582854
rect 363488 582586 363808 582618
rect 394208 583174 394528 583206
rect 394208 582938 394250 583174
rect 394486 582938 394528 583174
rect 394208 582854 394528 582938
rect 394208 582618 394250 582854
rect 394486 582618 394528 582854
rect 394208 582586 394528 582618
rect 424928 583174 425248 583206
rect 424928 582938 424970 583174
rect 425206 582938 425248 583174
rect 424928 582854 425248 582938
rect 424928 582618 424970 582854
rect 425206 582618 425248 582854
rect 424928 582586 425248 582618
rect 455648 583174 455968 583206
rect 455648 582938 455690 583174
rect 455926 582938 455968 583174
rect 455648 582854 455968 582938
rect 455648 582618 455690 582854
rect 455926 582618 455968 582854
rect 455648 582586 455968 582618
rect 486368 583174 486688 583206
rect 486368 582938 486410 583174
rect 486646 582938 486688 583174
rect 486368 582854 486688 582938
rect 486368 582618 486410 582854
rect 486646 582618 486688 582854
rect 486368 582586 486688 582618
rect 517088 583174 517408 583206
rect 517088 582938 517130 583174
rect 517366 582938 517408 583174
rect 517088 582854 517408 582938
rect 517088 582618 517130 582854
rect 517366 582618 517408 582854
rect 517088 582586 517408 582618
rect 547808 583174 548128 583206
rect 547808 582938 547850 583174
rect 548086 582938 548128 583174
rect 547808 582854 548128 582938
rect 547808 582618 547850 582854
rect 548086 582618 548128 582854
rect 547808 582586 548128 582618
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 10208 579454 10528 579486
rect 10208 579218 10250 579454
rect 10486 579218 10528 579454
rect 10208 579134 10528 579218
rect 10208 578898 10250 579134
rect 10486 578898 10528 579134
rect 10208 578866 10528 578898
rect 40928 579454 41248 579486
rect 40928 579218 40970 579454
rect 41206 579218 41248 579454
rect 40928 579134 41248 579218
rect 40928 578898 40970 579134
rect 41206 578898 41248 579134
rect 40928 578866 41248 578898
rect 71648 579454 71968 579486
rect 71648 579218 71690 579454
rect 71926 579218 71968 579454
rect 71648 579134 71968 579218
rect 71648 578898 71690 579134
rect 71926 578898 71968 579134
rect 71648 578866 71968 578898
rect 102368 579454 102688 579486
rect 102368 579218 102410 579454
rect 102646 579218 102688 579454
rect 102368 579134 102688 579218
rect 102368 578898 102410 579134
rect 102646 578898 102688 579134
rect 102368 578866 102688 578898
rect 133088 579454 133408 579486
rect 133088 579218 133130 579454
rect 133366 579218 133408 579454
rect 133088 579134 133408 579218
rect 133088 578898 133130 579134
rect 133366 578898 133408 579134
rect 133088 578866 133408 578898
rect 163808 579454 164128 579486
rect 163808 579218 163850 579454
rect 164086 579218 164128 579454
rect 163808 579134 164128 579218
rect 163808 578898 163850 579134
rect 164086 578898 164128 579134
rect 163808 578866 164128 578898
rect 194528 579454 194848 579486
rect 194528 579218 194570 579454
rect 194806 579218 194848 579454
rect 194528 579134 194848 579218
rect 194528 578898 194570 579134
rect 194806 578898 194848 579134
rect 194528 578866 194848 578898
rect 225248 579454 225568 579486
rect 225248 579218 225290 579454
rect 225526 579218 225568 579454
rect 225248 579134 225568 579218
rect 225248 578898 225290 579134
rect 225526 578898 225568 579134
rect 225248 578866 225568 578898
rect 255968 579454 256288 579486
rect 255968 579218 256010 579454
rect 256246 579218 256288 579454
rect 255968 579134 256288 579218
rect 255968 578898 256010 579134
rect 256246 578898 256288 579134
rect 255968 578866 256288 578898
rect 286688 579454 287008 579486
rect 286688 579218 286730 579454
rect 286966 579218 287008 579454
rect 286688 579134 287008 579218
rect 286688 578898 286730 579134
rect 286966 578898 287008 579134
rect 286688 578866 287008 578898
rect 317408 579454 317728 579486
rect 317408 579218 317450 579454
rect 317686 579218 317728 579454
rect 317408 579134 317728 579218
rect 317408 578898 317450 579134
rect 317686 578898 317728 579134
rect 317408 578866 317728 578898
rect 348128 579454 348448 579486
rect 348128 579218 348170 579454
rect 348406 579218 348448 579454
rect 348128 579134 348448 579218
rect 348128 578898 348170 579134
rect 348406 578898 348448 579134
rect 348128 578866 348448 578898
rect 378848 579454 379168 579486
rect 378848 579218 378890 579454
rect 379126 579218 379168 579454
rect 378848 579134 379168 579218
rect 378848 578898 378890 579134
rect 379126 578898 379168 579134
rect 378848 578866 379168 578898
rect 409568 579454 409888 579486
rect 409568 579218 409610 579454
rect 409846 579218 409888 579454
rect 409568 579134 409888 579218
rect 409568 578898 409610 579134
rect 409846 578898 409888 579134
rect 409568 578866 409888 578898
rect 440288 579454 440608 579486
rect 440288 579218 440330 579454
rect 440566 579218 440608 579454
rect 440288 579134 440608 579218
rect 440288 578898 440330 579134
rect 440566 578898 440608 579134
rect 440288 578866 440608 578898
rect 471008 579454 471328 579486
rect 471008 579218 471050 579454
rect 471286 579218 471328 579454
rect 471008 579134 471328 579218
rect 471008 578898 471050 579134
rect 471286 578898 471328 579134
rect 471008 578866 471328 578898
rect 501728 579454 502048 579486
rect 501728 579218 501770 579454
rect 502006 579218 502048 579454
rect 501728 579134 502048 579218
rect 501728 578898 501770 579134
rect 502006 578898 502048 579134
rect 501728 578866 502048 578898
rect 532448 579454 532768 579486
rect 532448 579218 532490 579454
rect 532726 579218 532768 579454
rect 532448 579134 532768 579218
rect 532448 578898 532490 579134
rect 532726 578898 532768 579134
rect 532448 578866 532768 578898
rect 563168 579454 563488 579486
rect 563168 579218 563210 579454
rect 563446 579218 563488 579454
rect 563168 579134 563488 579218
rect 563168 578898 563210 579134
rect 563446 578898 563488 579134
rect 563168 578866 563488 578898
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 25568 547174 25888 547206
rect 25568 546938 25610 547174
rect 25846 546938 25888 547174
rect 25568 546854 25888 546938
rect 25568 546618 25610 546854
rect 25846 546618 25888 546854
rect 25568 546586 25888 546618
rect 56288 547174 56608 547206
rect 56288 546938 56330 547174
rect 56566 546938 56608 547174
rect 56288 546854 56608 546938
rect 56288 546618 56330 546854
rect 56566 546618 56608 546854
rect 56288 546586 56608 546618
rect 87008 547174 87328 547206
rect 87008 546938 87050 547174
rect 87286 546938 87328 547174
rect 87008 546854 87328 546938
rect 87008 546618 87050 546854
rect 87286 546618 87328 546854
rect 87008 546586 87328 546618
rect 117728 547174 118048 547206
rect 117728 546938 117770 547174
rect 118006 546938 118048 547174
rect 117728 546854 118048 546938
rect 117728 546618 117770 546854
rect 118006 546618 118048 546854
rect 117728 546586 118048 546618
rect 148448 547174 148768 547206
rect 148448 546938 148490 547174
rect 148726 546938 148768 547174
rect 148448 546854 148768 546938
rect 148448 546618 148490 546854
rect 148726 546618 148768 546854
rect 148448 546586 148768 546618
rect 179168 547174 179488 547206
rect 179168 546938 179210 547174
rect 179446 546938 179488 547174
rect 179168 546854 179488 546938
rect 179168 546618 179210 546854
rect 179446 546618 179488 546854
rect 179168 546586 179488 546618
rect 209888 547174 210208 547206
rect 209888 546938 209930 547174
rect 210166 546938 210208 547174
rect 209888 546854 210208 546938
rect 209888 546618 209930 546854
rect 210166 546618 210208 546854
rect 209888 546586 210208 546618
rect 240608 547174 240928 547206
rect 240608 546938 240650 547174
rect 240886 546938 240928 547174
rect 240608 546854 240928 546938
rect 240608 546618 240650 546854
rect 240886 546618 240928 546854
rect 240608 546586 240928 546618
rect 271328 547174 271648 547206
rect 271328 546938 271370 547174
rect 271606 546938 271648 547174
rect 271328 546854 271648 546938
rect 271328 546618 271370 546854
rect 271606 546618 271648 546854
rect 271328 546586 271648 546618
rect 302048 547174 302368 547206
rect 302048 546938 302090 547174
rect 302326 546938 302368 547174
rect 302048 546854 302368 546938
rect 302048 546618 302090 546854
rect 302326 546618 302368 546854
rect 302048 546586 302368 546618
rect 332768 547174 333088 547206
rect 332768 546938 332810 547174
rect 333046 546938 333088 547174
rect 332768 546854 333088 546938
rect 332768 546618 332810 546854
rect 333046 546618 333088 546854
rect 332768 546586 333088 546618
rect 363488 547174 363808 547206
rect 363488 546938 363530 547174
rect 363766 546938 363808 547174
rect 363488 546854 363808 546938
rect 363488 546618 363530 546854
rect 363766 546618 363808 546854
rect 363488 546586 363808 546618
rect 394208 547174 394528 547206
rect 394208 546938 394250 547174
rect 394486 546938 394528 547174
rect 394208 546854 394528 546938
rect 394208 546618 394250 546854
rect 394486 546618 394528 546854
rect 394208 546586 394528 546618
rect 424928 547174 425248 547206
rect 424928 546938 424970 547174
rect 425206 546938 425248 547174
rect 424928 546854 425248 546938
rect 424928 546618 424970 546854
rect 425206 546618 425248 546854
rect 424928 546586 425248 546618
rect 455648 547174 455968 547206
rect 455648 546938 455690 547174
rect 455926 546938 455968 547174
rect 455648 546854 455968 546938
rect 455648 546618 455690 546854
rect 455926 546618 455968 546854
rect 455648 546586 455968 546618
rect 486368 547174 486688 547206
rect 486368 546938 486410 547174
rect 486646 546938 486688 547174
rect 486368 546854 486688 546938
rect 486368 546618 486410 546854
rect 486646 546618 486688 546854
rect 486368 546586 486688 546618
rect 517088 547174 517408 547206
rect 517088 546938 517130 547174
rect 517366 546938 517408 547174
rect 517088 546854 517408 546938
rect 517088 546618 517130 546854
rect 517366 546618 517408 546854
rect 517088 546586 517408 546618
rect 547808 547174 548128 547206
rect 547808 546938 547850 547174
rect 548086 546938 548128 547174
rect 547808 546854 548128 546938
rect 547808 546618 547850 546854
rect 548086 546618 548128 546854
rect 547808 546586 548128 546618
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 10208 543454 10528 543486
rect 10208 543218 10250 543454
rect 10486 543218 10528 543454
rect 10208 543134 10528 543218
rect 10208 542898 10250 543134
rect 10486 542898 10528 543134
rect 10208 542866 10528 542898
rect 40928 543454 41248 543486
rect 40928 543218 40970 543454
rect 41206 543218 41248 543454
rect 40928 543134 41248 543218
rect 40928 542898 40970 543134
rect 41206 542898 41248 543134
rect 40928 542866 41248 542898
rect 71648 543454 71968 543486
rect 71648 543218 71690 543454
rect 71926 543218 71968 543454
rect 71648 543134 71968 543218
rect 71648 542898 71690 543134
rect 71926 542898 71968 543134
rect 71648 542866 71968 542898
rect 102368 543454 102688 543486
rect 102368 543218 102410 543454
rect 102646 543218 102688 543454
rect 102368 543134 102688 543218
rect 102368 542898 102410 543134
rect 102646 542898 102688 543134
rect 102368 542866 102688 542898
rect 133088 543454 133408 543486
rect 133088 543218 133130 543454
rect 133366 543218 133408 543454
rect 133088 543134 133408 543218
rect 133088 542898 133130 543134
rect 133366 542898 133408 543134
rect 133088 542866 133408 542898
rect 163808 543454 164128 543486
rect 163808 543218 163850 543454
rect 164086 543218 164128 543454
rect 163808 543134 164128 543218
rect 163808 542898 163850 543134
rect 164086 542898 164128 543134
rect 163808 542866 164128 542898
rect 194528 543454 194848 543486
rect 194528 543218 194570 543454
rect 194806 543218 194848 543454
rect 194528 543134 194848 543218
rect 194528 542898 194570 543134
rect 194806 542898 194848 543134
rect 194528 542866 194848 542898
rect 225248 543454 225568 543486
rect 225248 543218 225290 543454
rect 225526 543218 225568 543454
rect 225248 543134 225568 543218
rect 225248 542898 225290 543134
rect 225526 542898 225568 543134
rect 225248 542866 225568 542898
rect 255968 543454 256288 543486
rect 255968 543218 256010 543454
rect 256246 543218 256288 543454
rect 255968 543134 256288 543218
rect 255968 542898 256010 543134
rect 256246 542898 256288 543134
rect 255968 542866 256288 542898
rect 286688 543454 287008 543486
rect 286688 543218 286730 543454
rect 286966 543218 287008 543454
rect 286688 543134 287008 543218
rect 286688 542898 286730 543134
rect 286966 542898 287008 543134
rect 286688 542866 287008 542898
rect 317408 543454 317728 543486
rect 317408 543218 317450 543454
rect 317686 543218 317728 543454
rect 317408 543134 317728 543218
rect 317408 542898 317450 543134
rect 317686 542898 317728 543134
rect 317408 542866 317728 542898
rect 348128 543454 348448 543486
rect 348128 543218 348170 543454
rect 348406 543218 348448 543454
rect 348128 543134 348448 543218
rect 348128 542898 348170 543134
rect 348406 542898 348448 543134
rect 348128 542866 348448 542898
rect 378848 543454 379168 543486
rect 378848 543218 378890 543454
rect 379126 543218 379168 543454
rect 378848 543134 379168 543218
rect 378848 542898 378890 543134
rect 379126 542898 379168 543134
rect 378848 542866 379168 542898
rect 409568 543454 409888 543486
rect 409568 543218 409610 543454
rect 409846 543218 409888 543454
rect 409568 543134 409888 543218
rect 409568 542898 409610 543134
rect 409846 542898 409888 543134
rect 409568 542866 409888 542898
rect 440288 543454 440608 543486
rect 440288 543218 440330 543454
rect 440566 543218 440608 543454
rect 440288 543134 440608 543218
rect 440288 542898 440330 543134
rect 440566 542898 440608 543134
rect 440288 542866 440608 542898
rect 471008 543454 471328 543486
rect 471008 543218 471050 543454
rect 471286 543218 471328 543454
rect 471008 543134 471328 543218
rect 471008 542898 471050 543134
rect 471286 542898 471328 543134
rect 471008 542866 471328 542898
rect 501728 543454 502048 543486
rect 501728 543218 501770 543454
rect 502006 543218 502048 543454
rect 501728 543134 502048 543218
rect 501728 542898 501770 543134
rect 502006 542898 502048 543134
rect 501728 542866 502048 542898
rect 532448 543454 532768 543486
rect 532448 543218 532490 543454
rect 532726 543218 532768 543454
rect 532448 543134 532768 543218
rect 532448 542898 532490 543134
rect 532726 542898 532768 543134
rect 532448 542866 532768 542898
rect 563168 543454 563488 543486
rect 563168 543218 563210 543454
rect 563446 543218 563488 543454
rect 563168 543134 563488 543218
rect 563168 542898 563210 543134
rect 563446 542898 563488 543134
rect 563168 542866 563488 542898
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 25568 511174 25888 511206
rect 25568 510938 25610 511174
rect 25846 510938 25888 511174
rect 25568 510854 25888 510938
rect 25568 510618 25610 510854
rect 25846 510618 25888 510854
rect 25568 510586 25888 510618
rect 56288 511174 56608 511206
rect 56288 510938 56330 511174
rect 56566 510938 56608 511174
rect 56288 510854 56608 510938
rect 56288 510618 56330 510854
rect 56566 510618 56608 510854
rect 56288 510586 56608 510618
rect 87008 511174 87328 511206
rect 87008 510938 87050 511174
rect 87286 510938 87328 511174
rect 87008 510854 87328 510938
rect 87008 510618 87050 510854
rect 87286 510618 87328 510854
rect 87008 510586 87328 510618
rect 117728 511174 118048 511206
rect 117728 510938 117770 511174
rect 118006 510938 118048 511174
rect 117728 510854 118048 510938
rect 117728 510618 117770 510854
rect 118006 510618 118048 510854
rect 117728 510586 118048 510618
rect 148448 511174 148768 511206
rect 148448 510938 148490 511174
rect 148726 510938 148768 511174
rect 148448 510854 148768 510938
rect 148448 510618 148490 510854
rect 148726 510618 148768 510854
rect 148448 510586 148768 510618
rect 179168 511174 179488 511206
rect 179168 510938 179210 511174
rect 179446 510938 179488 511174
rect 179168 510854 179488 510938
rect 179168 510618 179210 510854
rect 179446 510618 179488 510854
rect 179168 510586 179488 510618
rect 209888 511174 210208 511206
rect 209888 510938 209930 511174
rect 210166 510938 210208 511174
rect 209888 510854 210208 510938
rect 209888 510618 209930 510854
rect 210166 510618 210208 510854
rect 209888 510586 210208 510618
rect 240608 511174 240928 511206
rect 240608 510938 240650 511174
rect 240886 510938 240928 511174
rect 240608 510854 240928 510938
rect 240608 510618 240650 510854
rect 240886 510618 240928 510854
rect 240608 510586 240928 510618
rect 271328 511174 271648 511206
rect 271328 510938 271370 511174
rect 271606 510938 271648 511174
rect 271328 510854 271648 510938
rect 271328 510618 271370 510854
rect 271606 510618 271648 510854
rect 271328 510586 271648 510618
rect 302048 511174 302368 511206
rect 302048 510938 302090 511174
rect 302326 510938 302368 511174
rect 302048 510854 302368 510938
rect 302048 510618 302090 510854
rect 302326 510618 302368 510854
rect 302048 510586 302368 510618
rect 332768 511174 333088 511206
rect 332768 510938 332810 511174
rect 333046 510938 333088 511174
rect 332768 510854 333088 510938
rect 332768 510618 332810 510854
rect 333046 510618 333088 510854
rect 332768 510586 333088 510618
rect 363488 511174 363808 511206
rect 363488 510938 363530 511174
rect 363766 510938 363808 511174
rect 363488 510854 363808 510938
rect 363488 510618 363530 510854
rect 363766 510618 363808 510854
rect 363488 510586 363808 510618
rect 394208 511174 394528 511206
rect 394208 510938 394250 511174
rect 394486 510938 394528 511174
rect 394208 510854 394528 510938
rect 394208 510618 394250 510854
rect 394486 510618 394528 510854
rect 394208 510586 394528 510618
rect 424928 511174 425248 511206
rect 424928 510938 424970 511174
rect 425206 510938 425248 511174
rect 424928 510854 425248 510938
rect 424928 510618 424970 510854
rect 425206 510618 425248 510854
rect 424928 510586 425248 510618
rect 455648 511174 455968 511206
rect 455648 510938 455690 511174
rect 455926 510938 455968 511174
rect 455648 510854 455968 510938
rect 455648 510618 455690 510854
rect 455926 510618 455968 510854
rect 455648 510586 455968 510618
rect 486368 511174 486688 511206
rect 486368 510938 486410 511174
rect 486646 510938 486688 511174
rect 486368 510854 486688 510938
rect 486368 510618 486410 510854
rect 486646 510618 486688 510854
rect 486368 510586 486688 510618
rect 517088 511174 517408 511206
rect 517088 510938 517130 511174
rect 517366 510938 517408 511174
rect 517088 510854 517408 510938
rect 517088 510618 517130 510854
rect 517366 510618 517408 510854
rect 517088 510586 517408 510618
rect 547808 511174 548128 511206
rect 547808 510938 547850 511174
rect 548086 510938 548128 511174
rect 547808 510854 548128 510938
rect 547808 510618 547850 510854
rect 548086 510618 548128 510854
rect 547808 510586 548128 510618
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 10208 507454 10528 507486
rect 10208 507218 10250 507454
rect 10486 507218 10528 507454
rect 10208 507134 10528 507218
rect 10208 506898 10250 507134
rect 10486 506898 10528 507134
rect 10208 506866 10528 506898
rect 40928 507454 41248 507486
rect 40928 507218 40970 507454
rect 41206 507218 41248 507454
rect 40928 507134 41248 507218
rect 40928 506898 40970 507134
rect 41206 506898 41248 507134
rect 40928 506866 41248 506898
rect 71648 507454 71968 507486
rect 71648 507218 71690 507454
rect 71926 507218 71968 507454
rect 71648 507134 71968 507218
rect 71648 506898 71690 507134
rect 71926 506898 71968 507134
rect 71648 506866 71968 506898
rect 102368 507454 102688 507486
rect 102368 507218 102410 507454
rect 102646 507218 102688 507454
rect 102368 507134 102688 507218
rect 102368 506898 102410 507134
rect 102646 506898 102688 507134
rect 102368 506866 102688 506898
rect 133088 507454 133408 507486
rect 133088 507218 133130 507454
rect 133366 507218 133408 507454
rect 133088 507134 133408 507218
rect 133088 506898 133130 507134
rect 133366 506898 133408 507134
rect 133088 506866 133408 506898
rect 163808 507454 164128 507486
rect 163808 507218 163850 507454
rect 164086 507218 164128 507454
rect 163808 507134 164128 507218
rect 163808 506898 163850 507134
rect 164086 506898 164128 507134
rect 163808 506866 164128 506898
rect 194528 507454 194848 507486
rect 194528 507218 194570 507454
rect 194806 507218 194848 507454
rect 194528 507134 194848 507218
rect 194528 506898 194570 507134
rect 194806 506898 194848 507134
rect 194528 506866 194848 506898
rect 225248 507454 225568 507486
rect 225248 507218 225290 507454
rect 225526 507218 225568 507454
rect 225248 507134 225568 507218
rect 225248 506898 225290 507134
rect 225526 506898 225568 507134
rect 225248 506866 225568 506898
rect 255968 507454 256288 507486
rect 255968 507218 256010 507454
rect 256246 507218 256288 507454
rect 255968 507134 256288 507218
rect 255968 506898 256010 507134
rect 256246 506898 256288 507134
rect 255968 506866 256288 506898
rect 286688 507454 287008 507486
rect 286688 507218 286730 507454
rect 286966 507218 287008 507454
rect 286688 507134 287008 507218
rect 286688 506898 286730 507134
rect 286966 506898 287008 507134
rect 286688 506866 287008 506898
rect 317408 507454 317728 507486
rect 317408 507218 317450 507454
rect 317686 507218 317728 507454
rect 317408 507134 317728 507218
rect 317408 506898 317450 507134
rect 317686 506898 317728 507134
rect 317408 506866 317728 506898
rect 348128 507454 348448 507486
rect 348128 507218 348170 507454
rect 348406 507218 348448 507454
rect 348128 507134 348448 507218
rect 348128 506898 348170 507134
rect 348406 506898 348448 507134
rect 348128 506866 348448 506898
rect 378848 507454 379168 507486
rect 378848 507218 378890 507454
rect 379126 507218 379168 507454
rect 378848 507134 379168 507218
rect 378848 506898 378890 507134
rect 379126 506898 379168 507134
rect 378848 506866 379168 506898
rect 409568 507454 409888 507486
rect 409568 507218 409610 507454
rect 409846 507218 409888 507454
rect 409568 507134 409888 507218
rect 409568 506898 409610 507134
rect 409846 506898 409888 507134
rect 409568 506866 409888 506898
rect 440288 507454 440608 507486
rect 440288 507218 440330 507454
rect 440566 507218 440608 507454
rect 440288 507134 440608 507218
rect 440288 506898 440330 507134
rect 440566 506898 440608 507134
rect 440288 506866 440608 506898
rect 471008 507454 471328 507486
rect 471008 507218 471050 507454
rect 471286 507218 471328 507454
rect 471008 507134 471328 507218
rect 471008 506898 471050 507134
rect 471286 506898 471328 507134
rect 471008 506866 471328 506898
rect 501728 507454 502048 507486
rect 501728 507218 501770 507454
rect 502006 507218 502048 507454
rect 501728 507134 502048 507218
rect 501728 506898 501770 507134
rect 502006 506898 502048 507134
rect 501728 506866 502048 506898
rect 532448 507454 532768 507486
rect 532448 507218 532490 507454
rect 532726 507218 532768 507454
rect 532448 507134 532768 507218
rect 532448 506898 532490 507134
rect 532726 506898 532768 507134
rect 532448 506866 532768 506898
rect 563168 507454 563488 507486
rect 563168 507218 563210 507454
rect 563446 507218 563488 507454
rect 563168 507134 563488 507218
rect 563168 506898 563210 507134
rect 563446 506898 563488 507134
rect 563168 506866 563488 506898
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 25568 475174 25888 475206
rect 25568 474938 25610 475174
rect 25846 474938 25888 475174
rect 25568 474854 25888 474938
rect 25568 474618 25610 474854
rect 25846 474618 25888 474854
rect 25568 474586 25888 474618
rect 56288 475174 56608 475206
rect 56288 474938 56330 475174
rect 56566 474938 56608 475174
rect 56288 474854 56608 474938
rect 56288 474618 56330 474854
rect 56566 474618 56608 474854
rect 56288 474586 56608 474618
rect 87008 475174 87328 475206
rect 87008 474938 87050 475174
rect 87286 474938 87328 475174
rect 87008 474854 87328 474938
rect 87008 474618 87050 474854
rect 87286 474618 87328 474854
rect 87008 474586 87328 474618
rect 117728 475174 118048 475206
rect 117728 474938 117770 475174
rect 118006 474938 118048 475174
rect 117728 474854 118048 474938
rect 117728 474618 117770 474854
rect 118006 474618 118048 474854
rect 117728 474586 118048 474618
rect 148448 475174 148768 475206
rect 148448 474938 148490 475174
rect 148726 474938 148768 475174
rect 148448 474854 148768 474938
rect 148448 474618 148490 474854
rect 148726 474618 148768 474854
rect 148448 474586 148768 474618
rect 179168 475174 179488 475206
rect 179168 474938 179210 475174
rect 179446 474938 179488 475174
rect 179168 474854 179488 474938
rect 179168 474618 179210 474854
rect 179446 474618 179488 474854
rect 179168 474586 179488 474618
rect 209888 475174 210208 475206
rect 209888 474938 209930 475174
rect 210166 474938 210208 475174
rect 209888 474854 210208 474938
rect 209888 474618 209930 474854
rect 210166 474618 210208 474854
rect 209888 474586 210208 474618
rect 240608 475174 240928 475206
rect 240608 474938 240650 475174
rect 240886 474938 240928 475174
rect 240608 474854 240928 474938
rect 240608 474618 240650 474854
rect 240886 474618 240928 474854
rect 240608 474586 240928 474618
rect 271328 475174 271648 475206
rect 271328 474938 271370 475174
rect 271606 474938 271648 475174
rect 271328 474854 271648 474938
rect 271328 474618 271370 474854
rect 271606 474618 271648 474854
rect 271328 474586 271648 474618
rect 302048 475174 302368 475206
rect 302048 474938 302090 475174
rect 302326 474938 302368 475174
rect 302048 474854 302368 474938
rect 302048 474618 302090 474854
rect 302326 474618 302368 474854
rect 302048 474586 302368 474618
rect 332768 475174 333088 475206
rect 332768 474938 332810 475174
rect 333046 474938 333088 475174
rect 332768 474854 333088 474938
rect 332768 474618 332810 474854
rect 333046 474618 333088 474854
rect 332768 474586 333088 474618
rect 363488 475174 363808 475206
rect 363488 474938 363530 475174
rect 363766 474938 363808 475174
rect 363488 474854 363808 474938
rect 363488 474618 363530 474854
rect 363766 474618 363808 474854
rect 363488 474586 363808 474618
rect 394208 475174 394528 475206
rect 394208 474938 394250 475174
rect 394486 474938 394528 475174
rect 394208 474854 394528 474938
rect 394208 474618 394250 474854
rect 394486 474618 394528 474854
rect 394208 474586 394528 474618
rect 424928 475174 425248 475206
rect 424928 474938 424970 475174
rect 425206 474938 425248 475174
rect 424928 474854 425248 474938
rect 424928 474618 424970 474854
rect 425206 474618 425248 474854
rect 424928 474586 425248 474618
rect 455648 475174 455968 475206
rect 455648 474938 455690 475174
rect 455926 474938 455968 475174
rect 455648 474854 455968 474938
rect 455648 474618 455690 474854
rect 455926 474618 455968 474854
rect 455648 474586 455968 474618
rect 486368 475174 486688 475206
rect 486368 474938 486410 475174
rect 486646 474938 486688 475174
rect 486368 474854 486688 474938
rect 486368 474618 486410 474854
rect 486646 474618 486688 474854
rect 486368 474586 486688 474618
rect 517088 475174 517408 475206
rect 517088 474938 517130 475174
rect 517366 474938 517408 475174
rect 517088 474854 517408 474938
rect 517088 474618 517130 474854
rect 517366 474618 517408 474854
rect 517088 474586 517408 474618
rect 547808 475174 548128 475206
rect 547808 474938 547850 475174
rect 548086 474938 548128 475174
rect 547808 474854 548128 474938
rect 547808 474618 547850 474854
rect 548086 474618 548128 474854
rect 547808 474586 548128 474618
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 10208 471454 10528 471486
rect 10208 471218 10250 471454
rect 10486 471218 10528 471454
rect 10208 471134 10528 471218
rect 10208 470898 10250 471134
rect 10486 470898 10528 471134
rect 10208 470866 10528 470898
rect 40928 471454 41248 471486
rect 40928 471218 40970 471454
rect 41206 471218 41248 471454
rect 40928 471134 41248 471218
rect 40928 470898 40970 471134
rect 41206 470898 41248 471134
rect 40928 470866 41248 470898
rect 71648 471454 71968 471486
rect 71648 471218 71690 471454
rect 71926 471218 71968 471454
rect 71648 471134 71968 471218
rect 71648 470898 71690 471134
rect 71926 470898 71968 471134
rect 71648 470866 71968 470898
rect 102368 471454 102688 471486
rect 102368 471218 102410 471454
rect 102646 471218 102688 471454
rect 102368 471134 102688 471218
rect 102368 470898 102410 471134
rect 102646 470898 102688 471134
rect 102368 470866 102688 470898
rect 133088 471454 133408 471486
rect 133088 471218 133130 471454
rect 133366 471218 133408 471454
rect 133088 471134 133408 471218
rect 133088 470898 133130 471134
rect 133366 470898 133408 471134
rect 133088 470866 133408 470898
rect 163808 471454 164128 471486
rect 163808 471218 163850 471454
rect 164086 471218 164128 471454
rect 163808 471134 164128 471218
rect 163808 470898 163850 471134
rect 164086 470898 164128 471134
rect 163808 470866 164128 470898
rect 194528 471454 194848 471486
rect 194528 471218 194570 471454
rect 194806 471218 194848 471454
rect 194528 471134 194848 471218
rect 194528 470898 194570 471134
rect 194806 470898 194848 471134
rect 194528 470866 194848 470898
rect 225248 471454 225568 471486
rect 225248 471218 225290 471454
rect 225526 471218 225568 471454
rect 225248 471134 225568 471218
rect 225248 470898 225290 471134
rect 225526 470898 225568 471134
rect 225248 470866 225568 470898
rect 255968 471454 256288 471486
rect 255968 471218 256010 471454
rect 256246 471218 256288 471454
rect 255968 471134 256288 471218
rect 255968 470898 256010 471134
rect 256246 470898 256288 471134
rect 255968 470866 256288 470898
rect 286688 471454 287008 471486
rect 286688 471218 286730 471454
rect 286966 471218 287008 471454
rect 286688 471134 287008 471218
rect 286688 470898 286730 471134
rect 286966 470898 287008 471134
rect 286688 470866 287008 470898
rect 317408 471454 317728 471486
rect 317408 471218 317450 471454
rect 317686 471218 317728 471454
rect 317408 471134 317728 471218
rect 317408 470898 317450 471134
rect 317686 470898 317728 471134
rect 317408 470866 317728 470898
rect 348128 471454 348448 471486
rect 348128 471218 348170 471454
rect 348406 471218 348448 471454
rect 348128 471134 348448 471218
rect 348128 470898 348170 471134
rect 348406 470898 348448 471134
rect 348128 470866 348448 470898
rect 378848 471454 379168 471486
rect 378848 471218 378890 471454
rect 379126 471218 379168 471454
rect 378848 471134 379168 471218
rect 378848 470898 378890 471134
rect 379126 470898 379168 471134
rect 378848 470866 379168 470898
rect 409568 471454 409888 471486
rect 409568 471218 409610 471454
rect 409846 471218 409888 471454
rect 409568 471134 409888 471218
rect 409568 470898 409610 471134
rect 409846 470898 409888 471134
rect 409568 470866 409888 470898
rect 440288 471454 440608 471486
rect 440288 471218 440330 471454
rect 440566 471218 440608 471454
rect 440288 471134 440608 471218
rect 440288 470898 440330 471134
rect 440566 470898 440608 471134
rect 440288 470866 440608 470898
rect 471008 471454 471328 471486
rect 471008 471218 471050 471454
rect 471286 471218 471328 471454
rect 471008 471134 471328 471218
rect 471008 470898 471050 471134
rect 471286 470898 471328 471134
rect 471008 470866 471328 470898
rect 501728 471454 502048 471486
rect 501728 471218 501770 471454
rect 502006 471218 502048 471454
rect 501728 471134 502048 471218
rect 501728 470898 501770 471134
rect 502006 470898 502048 471134
rect 501728 470866 502048 470898
rect 532448 471454 532768 471486
rect 532448 471218 532490 471454
rect 532726 471218 532768 471454
rect 532448 471134 532768 471218
rect 532448 470898 532490 471134
rect 532726 470898 532768 471134
rect 532448 470866 532768 470898
rect 563168 471454 563488 471486
rect 563168 471218 563210 471454
rect 563446 471218 563488 471454
rect 563168 471134 563488 471218
rect 563168 470898 563210 471134
rect 563446 470898 563488 471134
rect 563168 470866 563488 470898
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 25568 439174 25888 439206
rect 25568 438938 25610 439174
rect 25846 438938 25888 439174
rect 25568 438854 25888 438938
rect 25568 438618 25610 438854
rect 25846 438618 25888 438854
rect 25568 438586 25888 438618
rect 56288 439174 56608 439206
rect 56288 438938 56330 439174
rect 56566 438938 56608 439174
rect 56288 438854 56608 438938
rect 56288 438618 56330 438854
rect 56566 438618 56608 438854
rect 56288 438586 56608 438618
rect 87008 439174 87328 439206
rect 87008 438938 87050 439174
rect 87286 438938 87328 439174
rect 87008 438854 87328 438938
rect 87008 438618 87050 438854
rect 87286 438618 87328 438854
rect 87008 438586 87328 438618
rect 117728 439174 118048 439206
rect 117728 438938 117770 439174
rect 118006 438938 118048 439174
rect 117728 438854 118048 438938
rect 117728 438618 117770 438854
rect 118006 438618 118048 438854
rect 117728 438586 118048 438618
rect 148448 439174 148768 439206
rect 148448 438938 148490 439174
rect 148726 438938 148768 439174
rect 148448 438854 148768 438938
rect 148448 438618 148490 438854
rect 148726 438618 148768 438854
rect 148448 438586 148768 438618
rect 179168 439174 179488 439206
rect 179168 438938 179210 439174
rect 179446 438938 179488 439174
rect 179168 438854 179488 438938
rect 179168 438618 179210 438854
rect 179446 438618 179488 438854
rect 179168 438586 179488 438618
rect 209888 439174 210208 439206
rect 209888 438938 209930 439174
rect 210166 438938 210208 439174
rect 209888 438854 210208 438938
rect 209888 438618 209930 438854
rect 210166 438618 210208 438854
rect 209888 438586 210208 438618
rect 240608 439174 240928 439206
rect 240608 438938 240650 439174
rect 240886 438938 240928 439174
rect 240608 438854 240928 438938
rect 240608 438618 240650 438854
rect 240886 438618 240928 438854
rect 240608 438586 240928 438618
rect 271328 439174 271648 439206
rect 271328 438938 271370 439174
rect 271606 438938 271648 439174
rect 271328 438854 271648 438938
rect 271328 438618 271370 438854
rect 271606 438618 271648 438854
rect 271328 438586 271648 438618
rect 302048 439174 302368 439206
rect 302048 438938 302090 439174
rect 302326 438938 302368 439174
rect 302048 438854 302368 438938
rect 302048 438618 302090 438854
rect 302326 438618 302368 438854
rect 302048 438586 302368 438618
rect 332768 439174 333088 439206
rect 332768 438938 332810 439174
rect 333046 438938 333088 439174
rect 332768 438854 333088 438938
rect 332768 438618 332810 438854
rect 333046 438618 333088 438854
rect 332768 438586 333088 438618
rect 363488 439174 363808 439206
rect 363488 438938 363530 439174
rect 363766 438938 363808 439174
rect 363488 438854 363808 438938
rect 363488 438618 363530 438854
rect 363766 438618 363808 438854
rect 363488 438586 363808 438618
rect 394208 439174 394528 439206
rect 394208 438938 394250 439174
rect 394486 438938 394528 439174
rect 394208 438854 394528 438938
rect 394208 438618 394250 438854
rect 394486 438618 394528 438854
rect 394208 438586 394528 438618
rect 424928 439174 425248 439206
rect 424928 438938 424970 439174
rect 425206 438938 425248 439174
rect 424928 438854 425248 438938
rect 424928 438618 424970 438854
rect 425206 438618 425248 438854
rect 424928 438586 425248 438618
rect 455648 439174 455968 439206
rect 455648 438938 455690 439174
rect 455926 438938 455968 439174
rect 455648 438854 455968 438938
rect 455648 438618 455690 438854
rect 455926 438618 455968 438854
rect 455648 438586 455968 438618
rect 486368 439174 486688 439206
rect 486368 438938 486410 439174
rect 486646 438938 486688 439174
rect 486368 438854 486688 438938
rect 486368 438618 486410 438854
rect 486646 438618 486688 438854
rect 486368 438586 486688 438618
rect 517088 439174 517408 439206
rect 517088 438938 517130 439174
rect 517366 438938 517408 439174
rect 517088 438854 517408 438938
rect 517088 438618 517130 438854
rect 517366 438618 517408 438854
rect 517088 438586 517408 438618
rect 547808 439174 548128 439206
rect 547808 438938 547850 439174
rect 548086 438938 548128 439174
rect 547808 438854 548128 438938
rect 547808 438618 547850 438854
rect 548086 438618 548128 438854
rect 547808 438586 548128 438618
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 10208 435454 10528 435486
rect 10208 435218 10250 435454
rect 10486 435218 10528 435454
rect 10208 435134 10528 435218
rect 10208 434898 10250 435134
rect 10486 434898 10528 435134
rect 10208 434866 10528 434898
rect 40928 435454 41248 435486
rect 40928 435218 40970 435454
rect 41206 435218 41248 435454
rect 40928 435134 41248 435218
rect 40928 434898 40970 435134
rect 41206 434898 41248 435134
rect 40928 434866 41248 434898
rect 71648 435454 71968 435486
rect 71648 435218 71690 435454
rect 71926 435218 71968 435454
rect 71648 435134 71968 435218
rect 71648 434898 71690 435134
rect 71926 434898 71968 435134
rect 71648 434866 71968 434898
rect 102368 435454 102688 435486
rect 102368 435218 102410 435454
rect 102646 435218 102688 435454
rect 102368 435134 102688 435218
rect 102368 434898 102410 435134
rect 102646 434898 102688 435134
rect 102368 434866 102688 434898
rect 133088 435454 133408 435486
rect 133088 435218 133130 435454
rect 133366 435218 133408 435454
rect 133088 435134 133408 435218
rect 133088 434898 133130 435134
rect 133366 434898 133408 435134
rect 133088 434866 133408 434898
rect 163808 435454 164128 435486
rect 163808 435218 163850 435454
rect 164086 435218 164128 435454
rect 163808 435134 164128 435218
rect 163808 434898 163850 435134
rect 164086 434898 164128 435134
rect 163808 434866 164128 434898
rect 194528 435454 194848 435486
rect 194528 435218 194570 435454
rect 194806 435218 194848 435454
rect 194528 435134 194848 435218
rect 194528 434898 194570 435134
rect 194806 434898 194848 435134
rect 194528 434866 194848 434898
rect 225248 435454 225568 435486
rect 225248 435218 225290 435454
rect 225526 435218 225568 435454
rect 225248 435134 225568 435218
rect 225248 434898 225290 435134
rect 225526 434898 225568 435134
rect 225248 434866 225568 434898
rect 255968 435454 256288 435486
rect 255968 435218 256010 435454
rect 256246 435218 256288 435454
rect 255968 435134 256288 435218
rect 255968 434898 256010 435134
rect 256246 434898 256288 435134
rect 255968 434866 256288 434898
rect 286688 435454 287008 435486
rect 286688 435218 286730 435454
rect 286966 435218 287008 435454
rect 286688 435134 287008 435218
rect 286688 434898 286730 435134
rect 286966 434898 287008 435134
rect 286688 434866 287008 434898
rect 317408 435454 317728 435486
rect 317408 435218 317450 435454
rect 317686 435218 317728 435454
rect 317408 435134 317728 435218
rect 317408 434898 317450 435134
rect 317686 434898 317728 435134
rect 317408 434866 317728 434898
rect 348128 435454 348448 435486
rect 348128 435218 348170 435454
rect 348406 435218 348448 435454
rect 348128 435134 348448 435218
rect 348128 434898 348170 435134
rect 348406 434898 348448 435134
rect 348128 434866 348448 434898
rect 378848 435454 379168 435486
rect 378848 435218 378890 435454
rect 379126 435218 379168 435454
rect 378848 435134 379168 435218
rect 378848 434898 378890 435134
rect 379126 434898 379168 435134
rect 378848 434866 379168 434898
rect 409568 435454 409888 435486
rect 409568 435218 409610 435454
rect 409846 435218 409888 435454
rect 409568 435134 409888 435218
rect 409568 434898 409610 435134
rect 409846 434898 409888 435134
rect 409568 434866 409888 434898
rect 440288 435454 440608 435486
rect 440288 435218 440330 435454
rect 440566 435218 440608 435454
rect 440288 435134 440608 435218
rect 440288 434898 440330 435134
rect 440566 434898 440608 435134
rect 440288 434866 440608 434898
rect 471008 435454 471328 435486
rect 471008 435218 471050 435454
rect 471286 435218 471328 435454
rect 471008 435134 471328 435218
rect 471008 434898 471050 435134
rect 471286 434898 471328 435134
rect 471008 434866 471328 434898
rect 501728 435454 502048 435486
rect 501728 435218 501770 435454
rect 502006 435218 502048 435454
rect 501728 435134 502048 435218
rect 501728 434898 501770 435134
rect 502006 434898 502048 435134
rect 501728 434866 502048 434898
rect 532448 435454 532768 435486
rect 532448 435218 532490 435454
rect 532726 435218 532768 435454
rect 532448 435134 532768 435218
rect 532448 434898 532490 435134
rect 532726 434898 532768 435134
rect 532448 434866 532768 434898
rect 563168 435454 563488 435486
rect 563168 435218 563210 435454
rect 563446 435218 563488 435454
rect 563168 435134 563488 435218
rect 563168 434898 563210 435134
rect 563446 434898 563488 435134
rect 563168 434866 563488 434898
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 25568 403174 25888 403206
rect 25568 402938 25610 403174
rect 25846 402938 25888 403174
rect 25568 402854 25888 402938
rect 25568 402618 25610 402854
rect 25846 402618 25888 402854
rect 25568 402586 25888 402618
rect 56288 403174 56608 403206
rect 56288 402938 56330 403174
rect 56566 402938 56608 403174
rect 56288 402854 56608 402938
rect 56288 402618 56330 402854
rect 56566 402618 56608 402854
rect 56288 402586 56608 402618
rect 87008 403174 87328 403206
rect 87008 402938 87050 403174
rect 87286 402938 87328 403174
rect 87008 402854 87328 402938
rect 87008 402618 87050 402854
rect 87286 402618 87328 402854
rect 87008 402586 87328 402618
rect 117728 403174 118048 403206
rect 117728 402938 117770 403174
rect 118006 402938 118048 403174
rect 117728 402854 118048 402938
rect 117728 402618 117770 402854
rect 118006 402618 118048 402854
rect 117728 402586 118048 402618
rect 148448 403174 148768 403206
rect 148448 402938 148490 403174
rect 148726 402938 148768 403174
rect 148448 402854 148768 402938
rect 148448 402618 148490 402854
rect 148726 402618 148768 402854
rect 148448 402586 148768 402618
rect 179168 403174 179488 403206
rect 179168 402938 179210 403174
rect 179446 402938 179488 403174
rect 179168 402854 179488 402938
rect 179168 402618 179210 402854
rect 179446 402618 179488 402854
rect 179168 402586 179488 402618
rect 209888 403174 210208 403206
rect 209888 402938 209930 403174
rect 210166 402938 210208 403174
rect 209888 402854 210208 402938
rect 209888 402618 209930 402854
rect 210166 402618 210208 402854
rect 209888 402586 210208 402618
rect 240608 403174 240928 403206
rect 240608 402938 240650 403174
rect 240886 402938 240928 403174
rect 240608 402854 240928 402938
rect 240608 402618 240650 402854
rect 240886 402618 240928 402854
rect 240608 402586 240928 402618
rect 271328 403174 271648 403206
rect 271328 402938 271370 403174
rect 271606 402938 271648 403174
rect 271328 402854 271648 402938
rect 271328 402618 271370 402854
rect 271606 402618 271648 402854
rect 271328 402586 271648 402618
rect 302048 403174 302368 403206
rect 302048 402938 302090 403174
rect 302326 402938 302368 403174
rect 302048 402854 302368 402938
rect 302048 402618 302090 402854
rect 302326 402618 302368 402854
rect 302048 402586 302368 402618
rect 332768 403174 333088 403206
rect 332768 402938 332810 403174
rect 333046 402938 333088 403174
rect 332768 402854 333088 402938
rect 332768 402618 332810 402854
rect 333046 402618 333088 402854
rect 332768 402586 333088 402618
rect 363488 403174 363808 403206
rect 363488 402938 363530 403174
rect 363766 402938 363808 403174
rect 363488 402854 363808 402938
rect 363488 402618 363530 402854
rect 363766 402618 363808 402854
rect 363488 402586 363808 402618
rect 394208 403174 394528 403206
rect 394208 402938 394250 403174
rect 394486 402938 394528 403174
rect 394208 402854 394528 402938
rect 394208 402618 394250 402854
rect 394486 402618 394528 402854
rect 394208 402586 394528 402618
rect 424928 403174 425248 403206
rect 424928 402938 424970 403174
rect 425206 402938 425248 403174
rect 424928 402854 425248 402938
rect 424928 402618 424970 402854
rect 425206 402618 425248 402854
rect 424928 402586 425248 402618
rect 455648 403174 455968 403206
rect 455648 402938 455690 403174
rect 455926 402938 455968 403174
rect 455648 402854 455968 402938
rect 455648 402618 455690 402854
rect 455926 402618 455968 402854
rect 455648 402586 455968 402618
rect 486368 403174 486688 403206
rect 486368 402938 486410 403174
rect 486646 402938 486688 403174
rect 486368 402854 486688 402938
rect 486368 402618 486410 402854
rect 486646 402618 486688 402854
rect 486368 402586 486688 402618
rect 517088 403174 517408 403206
rect 517088 402938 517130 403174
rect 517366 402938 517408 403174
rect 517088 402854 517408 402938
rect 517088 402618 517130 402854
rect 517366 402618 517408 402854
rect 517088 402586 517408 402618
rect 547808 403174 548128 403206
rect 547808 402938 547850 403174
rect 548086 402938 548128 403174
rect 547808 402854 548128 402938
rect 547808 402618 547850 402854
rect 548086 402618 548128 402854
rect 547808 402586 548128 402618
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 10208 399454 10528 399486
rect 10208 399218 10250 399454
rect 10486 399218 10528 399454
rect 10208 399134 10528 399218
rect 10208 398898 10250 399134
rect 10486 398898 10528 399134
rect 10208 398866 10528 398898
rect 40928 399454 41248 399486
rect 40928 399218 40970 399454
rect 41206 399218 41248 399454
rect 40928 399134 41248 399218
rect 40928 398898 40970 399134
rect 41206 398898 41248 399134
rect 40928 398866 41248 398898
rect 71648 399454 71968 399486
rect 71648 399218 71690 399454
rect 71926 399218 71968 399454
rect 71648 399134 71968 399218
rect 71648 398898 71690 399134
rect 71926 398898 71968 399134
rect 71648 398866 71968 398898
rect 102368 399454 102688 399486
rect 102368 399218 102410 399454
rect 102646 399218 102688 399454
rect 102368 399134 102688 399218
rect 102368 398898 102410 399134
rect 102646 398898 102688 399134
rect 102368 398866 102688 398898
rect 133088 399454 133408 399486
rect 133088 399218 133130 399454
rect 133366 399218 133408 399454
rect 133088 399134 133408 399218
rect 133088 398898 133130 399134
rect 133366 398898 133408 399134
rect 133088 398866 133408 398898
rect 163808 399454 164128 399486
rect 163808 399218 163850 399454
rect 164086 399218 164128 399454
rect 163808 399134 164128 399218
rect 163808 398898 163850 399134
rect 164086 398898 164128 399134
rect 163808 398866 164128 398898
rect 194528 399454 194848 399486
rect 194528 399218 194570 399454
rect 194806 399218 194848 399454
rect 194528 399134 194848 399218
rect 194528 398898 194570 399134
rect 194806 398898 194848 399134
rect 194528 398866 194848 398898
rect 225248 399454 225568 399486
rect 225248 399218 225290 399454
rect 225526 399218 225568 399454
rect 225248 399134 225568 399218
rect 225248 398898 225290 399134
rect 225526 398898 225568 399134
rect 225248 398866 225568 398898
rect 255968 399454 256288 399486
rect 255968 399218 256010 399454
rect 256246 399218 256288 399454
rect 255968 399134 256288 399218
rect 255968 398898 256010 399134
rect 256246 398898 256288 399134
rect 255968 398866 256288 398898
rect 286688 399454 287008 399486
rect 286688 399218 286730 399454
rect 286966 399218 287008 399454
rect 286688 399134 287008 399218
rect 286688 398898 286730 399134
rect 286966 398898 287008 399134
rect 286688 398866 287008 398898
rect 317408 399454 317728 399486
rect 317408 399218 317450 399454
rect 317686 399218 317728 399454
rect 317408 399134 317728 399218
rect 317408 398898 317450 399134
rect 317686 398898 317728 399134
rect 317408 398866 317728 398898
rect 348128 399454 348448 399486
rect 348128 399218 348170 399454
rect 348406 399218 348448 399454
rect 348128 399134 348448 399218
rect 348128 398898 348170 399134
rect 348406 398898 348448 399134
rect 348128 398866 348448 398898
rect 378848 399454 379168 399486
rect 378848 399218 378890 399454
rect 379126 399218 379168 399454
rect 378848 399134 379168 399218
rect 378848 398898 378890 399134
rect 379126 398898 379168 399134
rect 378848 398866 379168 398898
rect 409568 399454 409888 399486
rect 409568 399218 409610 399454
rect 409846 399218 409888 399454
rect 409568 399134 409888 399218
rect 409568 398898 409610 399134
rect 409846 398898 409888 399134
rect 409568 398866 409888 398898
rect 440288 399454 440608 399486
rect 440288 399218 440330 399454
rect 440566 399218 440608 399454
rect 440288 399134 440608 399218
rect 440288 398898 440330 399134
rect 440566 398898 440608 399134
rect 440288 398866 440608 398898
rect 471008 399454 471328 399486
rect 471008 399218 471050 399454
rect 471286 399218 471328 399454
rect 471008 399134 471328 399218
rect 471008 398898 471050 399134
rect 471286 398898 471328 399134
rect 471008 398866 471328 398898
rect 501728 399454 502048 399486
rect 501728 399218 501770 399454
rect 502006 399218 502048 399454
rect 501728 399134 502048 399218
rect 501728 398898 501770 399134
rect 502006 398898 502048 399134
rect 501728 398866 502048 398898
rect 532448 399454 532768 399486
rect 532448 399218 532490 399454
rect 532726 399218 532768 399454
rect 532448 399134 532768 399218
rect 532448 398898 532490 399134
rect 532726 398898 532768 399134
rect 532448 398866 532768 398898
rect 563168 399454 563488 399486
rect 563168 399218 563210 399454
rect 563446 399218 563488 399454
rect 563168 399134 563488 399218
rect 563168 398898 563210 399134
rect 563446 398898 563488 399134
rect 563168 398866 563488 398898
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 25568 367174 25888 367206
rect 25568 366938 25610 367174
rect 25846 366938 25888 367174
rect 25568 366854 25888 366938
rect 25568 366618 25610 366854
rect 25846 366618 25888 366854
rect 25568 366586 25888 366618
rect 56288 367174 56608 367206
rect 56288 366938 56330 367174
rect 56566 366938 56608 367174
rect 56288 366854 56608 366938
rect 56288 366618 56330 366854
rect 56566 366618 56608 366854
rect 56288 366586 56608 366618
rect 87008 367174 87328 367206
rect 87008 366938 87050 367174
rect 87286 366938 87328 367174
rect 87008 366854 87328 366938
rect 87008 366618 87050 366854
rect 87286 366618 87328 366854
rect 87008 366586 87328 366618
rect 117728 367174 118048 367206
rect 117728 366938 117770 367174
rect 118006 366938 118048 367174
rect 117728 366854 118048 366938
rect 117728 366618 117770 366854
rect 118006 366618 118048 366854
rect 117728 366586 118048 366618
rect 148448 367174 148768 367206
rect 148448 366938 148490 367174
rect 148726 366938 148768 367174
rect 148448 366854 148768 366938
rect 148448 366618 148490 366854
rect 148726 366618 148768 366854
rect 148448 366586 148768 366618
rect 179168 367174 179488 367206
rect 179168 366938 179210 367174
rect 179446 366938 179488 367174
rect 179168 366854 179488 366938
rect 179168 366618 179210 366854
rect 179446 366618 179488 366854
rect 179168 366586 179488 366618
rect 209888 367174 210208 367206
rect 209888 366938 209930 367174
rect 210166 366938 210208 367174
rect 209888 366854 210208 366938
rect 209888 366618 209930 366854
rect 210166 366618 210208 366854
rect 209888 366586 210208 366618
rect 240608 367174 240928 367206
rect 240608 366938 240650 367174
rect 240886 366938 240928 367174
rect 240608 366854 240928 366938
rect 240608 366618 240650 366854
rect 240886 366618 240928 366854
rect 240608 366586 240928 366618
rect 271328 367174 271648 367206
rect 271328 366938 271370 367174
rect 271606 366938 271648 367174
rect 271328 366854 271648 366938
rect 271328 366618 271370 366854
rect 271606 366618 271648 366854
rect 271328 366586 271648 366618
rect 302048 367174 302368 367206
rect 302048 366938 302090 367174
rect 302326 366938 302368 367174
rect 302048 366854 302368 366938
rect 302048 366618 302090 366854
rect 302326 366618 302368 366854
rect 302048 366586 302368 366618
rect 332768 367174 333088 367206
rect 332768 366938 332810 367174
rect 333046 366938 333088 367174
rect 332768 366854 333088 366938
rect 332768 366618 332810 366854
rect 333046 366618 333088 366854
rect 332768 366586 333088 366618
rect 363488 367174 363808 367206
rect 363488 366938 363530 367174
rect 363766 366938 363808 367174
rect 363488 366854 363808 366938
rect 363488 366618 363530 366854
rect 363766 366618 363808 366854
rect 363488 366586 363808 366618
rect 394208 367174 394528 367206
rect 394208 366938 394250 367174
rect 394486 366938 394528 367174
rect 394208 366854 394528 366938
rect 394208 366618 394250 366854
rect 394486 366618 394528 366854
rect 394208 366586 394528 366618
rect 424928 367174 425248 367206
rect 424928 366938 424970 367174
rect 425206 366938 425248 367174
rect 424928 366854 425248 366938
rect 424928 366618 424970 366854
rect 425206 366618 425248 366854
rect 424928 366586 425248 366618
rect 455648 367174 455968 367206
rect 455648 366938 455690 367174
rect 455926 366938 455968 367174
rect 455648 366854 455968 366938
rect 455648 366618 455690 366854
rect 455926 366618 455968 366854
rect 455648 366586 455968 366618
rect 486368 367174 486688 367206
rect 486368 366938 486410 367174
rect 486646 366938 486688 367174
rect 486368 366854 486688 366938
rect 486368 366618 486410 366854
rect 486646 366618 486688 366854
rect 486368 366586 486688 366618
rect 517088 367174 517408 367206
rect 517088 366938 517130 367174
rect 517366 366938 517408 367174
rect 517088 366854 517408 366938
rect 517088 366618 517130 366854
rect 517366 366618 517408 366854
rect 517088 366586 517408 366618
rect 547808 367174 548128 367206
rect 547808 366938 547850 367174
rect 548086 366938 548128 367174
rect 547808 366854 548128 366938
rect 547808 366618 547850 366854
rect 548086 366618 548128 366854
rect 547808 366586 548128 366618
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 10208 363454 10528 363486
rect 10208 363218 10250 363454
rect 10486 363218 10528 363454
rect 10208 363134 10528 363218
rect 10208 362898 10250 363134
rect 10486 362898 10528 363134
rect 10208 362866 10528 362898
rect 40928 363454 41248 363486
rect 40928 363218 40970 363454
rect 41206 363218 41248 363454
rect 40928 363134 41248 363218
rect 40928 362898 40970 363134
rect 41206 362898 41248 363134
rect 40928 362866 41248 362898
rect 71648 363454 71968 363486
rect 71648 363218 71690 363454
rect 71926 363218 71968 363454
rect 71648 363134 71968 363218
rect 71648 362898 71690 363134
rect 71926 362898 71968 363134
rect 71648 362866 71968 362898
rect 102368 363454 102688 363486
rect 102368 363218 102410 363454
rect 102646 363218 102688 363454
rect 102368 363134 102688 363218
rect 102368 362898 102410 363134
rect 102646 362898 102688 363134
rect 102368 362866 102688 362898
rect 133088 363454 133408 363486
rect 133088 363218 133130 363454
rect 133366 363218 133408 363454
rect 133088 363134 133408 363218
rect 133088 362898 133130 363134
rect 133366 362898 133408 363134
rect 133088 362866 133408 362898
rect 163808 363454 164128 363486
rect 163808 363218 163850 363454
rect 164086 363218 164128 363454
rect 163808 363134 164128 363218
rect 163808 362898 163850 363134
rect 164086 362898 164128 363134
rect 163808 362866 164128 362898
rect 194528 363454 194848 363486
rect 194528 363218 194570 363454
rect 194806 363218 194848 363454
rect 194528 363134 194848 363218
rect 194528 362898 194570 363134
rect 194806 362898 194848 363134
rect 194528 362866 194848 362898
rect 225248 363454 225568 363486
rect 225248 363218 225290 363454
rect 225526 363218 225568 363454
rect 225248 363134 225568 363218
rect 225248 362898 225290 363134
rect 225526 362898 225568 363134
rect 225248 362866 225568 362898
rect 255968 363454 256288 363486
rect 255968 363218 256010 363454
rect 256246 363218 256288 363454
rect 255968 363134 256288 363218
rect 255968 362898 256010 363134
rect 256246 362898 256288 363134
rect 255968 362866 256288 362898
rect 286688 363454 287008 363486
rect 286688 363218 286730 363454
rect 286966 363218 287008 363454
rect 286688 363134 287008 363218
rect 286688 362898 286730 363134
rect 286966 362898 287008 363134
rect 286688 362866 287008 362898
rect 317408 363454 317728 363486
rect 317408 363218 317450 363454
rect 317686 363218 317728 363454
rect 317408 363134 317728 363218
rect 317408 362898 317450 363134
rect 317686 362898 317728 363134
rect 317408 362866 317728 362898
rect 348128 363454 348448 363486
rect 348128 363218 348170 363454
rect 348406 363218 348448 363454
rect 348128 363134 348448 363218
rect 348128 362898 348170 363134
rect 348406 362898 348448 363134
rect 348128 362866 348448 362898
rect 378848 363454 379168 363486
rect 378848 363218 378890 363454
rect 379126 363218 379168 363454
rect 378848 363134 379168 363218
rect 378848 362898 378890 363134
rect 379126 362898 379168 363134
rect 378848 362866 379168 362898
rect 409568 363454 409888 363486
rect 409568 363218 409610 363454
rect 409846 363218 409888 363454
rect 409568 363134 409888 363218
rect 409568 362898 409610 363134
rect 409846 362898 409888 363134
rect 409568 362866 409888 362898
rect 440288 363454 440608 363486
rect 440288 363218 440330 363454
rect 440566 363218 440608 363454
rect 440288 363134 440608 363218
rect 440288 362898 440330 363134
rect 440566 362898 440608 363134
rect 440288 362866 440608 362898
rect 471008 363454 471328 363486
rect 471008 363218 471050 363454
rect 471286 363218 471328 363454
rect 471008 363134 471328 363218
rect 471008 362898 471050 363134
rect 471286 362898 471328 363134
rect 471008 362866 471328 362898
rect 501728 363454 502048 363486
rect 501728 363218 501770 363454
rect 502006 363218 502048 363454
rect 501728 363134 502048 363218
rect 501728 362898 501770 363134
rect 502006 362898 502048 363134
rect 501728 362866 502048 362898
rect 532448 363454 532768 363486
rect 532448 363218 532490 363454
rect 532726 363218 532768 363454
rect 532448 363134 532768 363218
rect 532448 362898 532490 363134
rect 532726 362898 532768 363134
rect 532448 362866 532768 362898
rect 563168 363454 563488 363486
rect 563168 363218 563210 363454
rect 563446 363218 563488 363454
rect 563168 363134 563488 363218
rect 563168 362898 563210 363134
rect 563446 362898 563488 363134
rect 563168 362866 563488 362898
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 25568 331174 25888 331206
rect 25568 330938 25610 331174
rect 25846 330938 25888 331174
rect 25568 330854 25888 330938
rect 25568 330618 25610 330854
rect 25846 330618 25888 330854
rect 25568 330586 25888 330618
rect 56288 331174 56608 331206
rect 56288 330938 56330 331174
rect 56566 330938 56608 331174
rect 56288 330854 56608 330938
rect 56288 330618 56330 330854
rect 56566 330618 56608 330854
rect 56288 330586 56608 330618
rect 87008 331174 87328 331206
rect 87008 330938 87050 331174
rect 87286 330938 87328 331174
rect 87008 330854 87328 330938
rect 87008 330618 87050 330854
rect 87286 330618 87328 330854
rect 87008 330586 87328 330618
rect 117728 331174 118048 331206
rect 117728 330938 117770 331174
rect 118006 330938 118048 331174
rect 117728 330854 118048 330938
rect 117728 330618 117770 330854
rect 118006 330618 118048 330854
rect 117728 330586 118048 330618
rect 148448 331174 148768 331206
rect 148448 330938 148490 331174
rect 148726 330938 148768 331174
rect 148448 330854 148768 330938
rect 148448 330618 148490 330854
rect 148726 330618 148768 330854
rect 148448 330586 148768 330618
rect 179168 331174 179488 331206
rect 179168 330938 179210 331174
rect 179446 330938 179488 331174
rect 179168 330854 179488 330938
rect 179168 330618 179210 330854
rect 179446 330618 179488 330854
rect 179168 330586 179488 330618
rect 209888 331174 210208 331206
rect 209888 330938 209930 331174
rect 210166 330938 210208 331174
rect 209888 330854 210208 330938
rect 209888 330618 209930 330854
rect 210166 330618 210208 330854
rect 209888 330586 210208 330618
rect 240608 331174 240928 331206
rect 240608 330938 240650 331174
rect 240886 330938 240928 331174
rect 240608 330854 240928 330938
rect 240608 330618 240650 330854
rect 240886 330618 240928 330854
rect 240608 330586 240928 330618
rect 271328 331174 271648 331206
rect 271328 330938 271370 331174
rect 271606 330938 271648 331174
rect 271328 330854 271648 330938
rect 271328 330618 271370 330854
rect 271606 330618 271648 330854
rect 271328 330586 271648 330618
rect 302048 331174 302368 331206
rect 302048 330938 302090 331174
rect 302326 330938 302368 331174
rect 302048 330854 302368 330938
rect 302048 330618 302090 330854
rect 302326 330618 302368 330854
rect 302048 330586 302368 330618
rect 332768 331174 333088 331206
rect 332768 330938 332810 331174
rect 333046 330938 333088 331174
rect 332768 330854 333088 330938
rect 332768 330618 332810 330854
rect 333046 330618 333088 330854
rect 332768 330586 333088 330618
rect 363488 331174 363808 331206
rect 363488 330938 363530 331174
rect 363766 330938 363808 331174
rect 363488 330854 363808 330938
rect 363488 330618 363530 330854
rect 363766 330618 363808 330854
rect 363488 330586 363808 330618
rect 394208 331174 394528 331206
rect 394208 330938 394250 331174
rect 394486 330938 394528 331174
rect 394208 330854 394528 330938
rect 394208 330618 394250 330854
rect 394486 330618 394528 330854
rect 394208 330586 394528 330618
rect 424928 331174 425248 331206
rect 424928 330938 424970 331174
rect 425206 330938 425248 331174
rect 424928 330854 425248 330938
rect 424928 330618 424970 330854
rect 425206 330618 425248 330854
rect 424928 330586 425248 330618
rect 455648 331174 455968 331206
rect 455648 330938 455690 331174
rect 455926 330938 455968 331174
rect 455648 330854 455968 330938
rect 455648 330618 455690 330854
rect 455926 330618 455968 330854
rect 455648 330586 455968 330618
rect 486368 331174 486688 331206
rect 486368 330938 486410 331174
rect 486646 330938 486688 331174
rect 486368 330854 486688 330938
rect 486368 330618 486410 330854
rect 486646 330618 486688 330854
rect 486368 330586 486688 330618
rect 517088 331174 517408 331206
rect 517088 330938 517130 331174
rect 517366 330938 517408 331174
rect 517088 330854 517408 330938
rect 517088 330618 517130 330854
rect 517366 330618 517408 330854
rect 517088 330586 517408 330618
rect 547808 331174 548128 331206
rect 547808 330938 547850 331174
rect 548086 330938 548128 331174
rect 547808 330854 548128 330938
rect 547808 330618 547850 330854
rect 548086 330618 548128 330854
rect 547808 330586 548128 330618
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 10208 327454 10528 327486
rect 10208 327218 10250 327454
rect 10486 327218 10528 327454
rect 10208 327134 10528 327218
rect 10208 326898 10250 327134
rect 10486 326898 10528 327134
rect 10208 326866 10528 326898
rect 40928 327454 41248 327486
rect 40928 327218 40970 327454
rect 41206 327218 41248 327454
rect 40928 327134 41248 327218
rect 40928 326898 40970 327134
rect 41206 326898 41248 327134
rect 40928 326866 41248 326898
rect 71648 327454 71968 327486
rect 71648 327218 71690 327454
rect 71926 327218 71968 327454
rect 71648 327134 71968 327218
rect 71648 326898 71690 327134
rect 71926 326898 71968 327134
rect 71648 326866 71968 326898
rect 102368 327454 102688 327486
rect 102368 327218 102410 327454
rect 102646 327218 102688 327454
rect 102368 327134 102688 327218
rect 102368 326898 102410 327134
rect 102646 326898 102688 327134
rect 102368 326866 102688 326898
rect 133088 327454 133408 327486
rect 133088 327218 133130 327454
rect 133366 327218 133408 327454
rect 133088 327134 133408 327218
rect 133088 326898 133130 327134
rect 133366 326898 133408 327134
rect 133088 326866 133408 326898
rect 163808 327454 164128 327486
rect 163808 327218 163850 327454
rect 164086 327218 164128 327454
rect 163808 327134 164128 327218
rect 163808 326898 163850 327134
rect 164086 326898 164128 327134
rect 163808 326866 164128 326898
rect 194528 327454 194848 327486
rect 194528 327218 194570 327454
rect 194806 327218 194848 327454
rect 194528 327134 194848 327218
rect 194528 326898 194570 327134
rect 194806 326898 194848 327134
rect 194528 326866 194848 326898
rect 225248 327454 225568 327486
rect 225248 327218 225290 327454
rect 225526 327218 225568 327454
rect 225248 327134 225568 327218
rect 225248 326898 225290 327134
rect 225526 326898 225568 327134
rect 225248 326866 225568 326898
rect 255968 327454 256288 327486
rect 255968 327218 256010 327454
rect 256246 327218 256288 327454
rect 255968 327134 256288 327218
rect 255968 326898 256010 327134
rect 256246 326898 256288 327134
rect 255968 326866 256288 326898
rect 286688 327454 287008 327486
rect 286688 327218 286730 327454
rect 286966 327218 287008 327454
rect 286688 327134 287008 327218
rect 286688 326898 286730 327134
rect 286966 326898 287008 327134
rect 286688 326866 287008 326898
rect 317408 327454 317728 327486
rect 317408 327218 317450 327454
rect 317686 327218 317728 327454
rect 317408 327134 317728 327218
rect 317408 326898 317450 327134
rect 317686 326898 317728 327134
rect 317408 326866 317728 326898
rect 348128 327454 348448 327486
rect 348128 327218 348170 327454
rect 348406 327218 348448 327454
rect 348128 327134 348448 327218
rect 348128 326898 348170 327134
rect 348406 326898 348448 327134
rect 348128 326866 348448 326898
rect 378848 327454 379168 327486
rect 378848 327218 378890 327454
rect 379126 327218 379168 327454
rect 378848 327134 379168 327218
rect 378848 326898 378890 327134
rect 379126 326898 379168 327134
rect 378848 326866 379168 326898
rect 409568 327454 409888 327486
rect 409568 327218 409610 327454
rect 409846 327218 409888 327454
rect 409568 327134 409888 327218
rect 409568 326898 409610 327134
rect 409846 326898 409888 327134
rect 409568 326866 409888 326898
rect 440288 327454 440608 327486
rect 440288 327218 440330 327454
rect 440566 327218 440608 327454
rect 440288 327134 440608 327218
rect 440288 326898 440330 327134
rect 440566 326898 440608 327134
rect 440288 326866 440608 326898
rect 471008 327454 471328 327486
rect 471008 327218 471050 327454
rect 471286 327218 471328 327454
rect 471008 327134 471328 327218
rect 471008 326898 471050 327134
rect 471286 326898 471328 327134
rect 471008 326866 471328 326898
rect 501728 327454 502048 327486
rect 501728 327218 501770 327454
rect 502006 327218 502048 327454
rect 501728 327134 502048 327218
rect 501728 326898 501770 327134
rect 502006 326898 502048 327134
rect 501728 326866 502048 326898
rect 532448 327454 532768 327486
rect 532448 327218 532490 327454
rect 532726 327218 532768 327454
rect 532448 327134 532768 327218
rect 532448 326898 532490 327134
rect 532726 326898 532768 327134
rect 532448 326866 532768 326898
rect 563168 327454 563488 327486
rect 563168 327218 563210 327454
rect 563446 327218 563488 327454
rect 563168 327134 563488 327218
rect 563168 326898 563210 327134
rect 563446 326898 563488 327134
rect 563168 326866 563488 326898
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 25568 295174 25888 295206
rect 25568 294938 25610 295174
rect 25846 294938 25888 295174
rect 25568 294854 25888 294938
rect 25568 294618 25610 294854
rect 25846 294618 25888 294854
rect 25568 294586 25888 294618
rect 56288 295174 56608 295206
rect 56288 294938 56330 295174
rect 56566 294938 56608 295174
rect 56288 294854 56608 294938
rect 56288 294618 56330 294854
rect 56566 294618 56608 294854
rect 56288 294586 56608 294618
rect 87008 295174 87328 295206
rect 87008 294938 87050 295174
rect 87286 294938 87328 295174
rect 87008 294854 87328 294938
rect 87008 294618 87050 294854
rect 87286 294618 87328 294854
rect 87008 294586 87328 294618
rect 117728 295174 118048 295206
rect 117728 294938 117770 295174
rect 118006 294938 118048 295174
rect 117728 294854 118048 294938
rect 117728 294618 117770 294854
rect 118006 294618 118048 294854
rect 117728 294586 118048 294618
rect 148448 295174 148768 295206
rect 148448 294938 148490 295174
rect 148726 294938 148768 295174
rect 148448 294854 148768 294938
rect 148448 294618 148490 294854
rect 148726 294618 148768 294854
rect 148448 294586 148768 294618
rect 179168 295174 179488 295206
rect 179168 294938 179210 295174
rect 179446 294938 179488 295174
rect 179168 294854 179488 294938
rect 179168 294618 179210 294854
rect 179446 294618 179488 294854
rect 179168 294586 179488 294618
rect 209888 295174 210208 295206
rect 209888 294938 209930 295174
rect 210166 294938 210208 295174
rect 209888 294854 210208 294938
rect 209888 294618 209930 294854
rect 210166 294618 210208 294854
rect 209888 294586 210208 294618
rect 240608 295174 240928 295206
rect 240608 294938 240650 295174
rect 240886 294938 240928 295174
rect 240608 294854 240928 294938
rect 240608 294618 240650 294854
rect 240886 294618 240928 294854
rect 240608 294586 240928 294618
rect 271328 295174 271648 295206
rect 271328 294938 271370 295174
rect 271606 294938 271648 295174
rect 271328 294854 271648 294938
rect 271328 294618 271370 294854
rect 271606 294618 271648 294854
rect 271328 294586 271648 294618
rect 302048 295174 302368 295206
rect 302048 294938 302090 295174
rect 302326 294938 302368 295174
rect 302048 294854 302368 294938
rect 302048 294618 302090 294854
rect 302326 294618 302368 294854
rect 302048 294586 302368 294618
rect 332768 295174 333088 295206
rect 332768 294938 332810 295174
rect 333046 294938 333088 295174
rect 332768 294854 333088 294938
rect 332768 294618 332810 294854
rect 333046 294618 333088 294854
rect 332768 294586 333088 294618
rect 363488 295174 363808 295206
rect 363488 294938 363530 295174
rect 363766 294938 363808 295174
rect 363488 294854 363808 294938
rect 363488 294618 363530 294854
rect 363766 294618 363808 294854
rect 363488 294586 363808 294618
rect 394208 295174 394528 295206
rect 394208 294938 394250 295174
rect 394486 294938 394528 295174
rect 394208 294854 394528 294938
rect 394208 294618 394250 294854
rect 394486 294618 394528 294854
rect 394208 294586 394528 294618
rect 424928 295174 425248 295206
rect 424928 294938 424970 295174
rect 425206 294938 425248 295174
rect 424928 294854 425248 294938
rect 424928 294618 424970 294854
rect 425206 294618 425248 294854
rect 424928 294586 425248 294618
rect 455648 295174 455968 295206
rect 455648 294938 455690 295174
rect 455926 294938 455968 295174
rect 455648 294854 455968 294938
rect 455648 294618 455690 294854
rect 455926 294618 455968 294854
rect 455648 294586 455968 294618
rect 486368 295174 486688 295206
rect 486368 294938 486410 295174
rect 486646 294938 486688 295174
rect 486368 294854 486688 294938
rect 486368 294618 486410 294854
rect 486646 294618 486688 294854
rect 486368 294586 486688 294618
rect 517088 295174 517408 295206
rect 517088 294938 517130 295174
rect 517366 294938 517408 295174
rect 517088 294854 517408 294938
rect 517088 294618 517130 294854
rect 517366 294618 517408 294854
rect 517088 294586 517408 294618
rect 547808 295174 548128 295206
rect 547808 294938 547850 295174
rect 548086 294938 548128 295174
rect 547808 294854 548128 294938
rect 547808 294618 547850 294854
rect 548086 294618 548128 294854
rect 547808 294586 548128 294618
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 10208 291454 10528 291486
rect 10208 291218 10250 291454
rect 10486 291218 10528 291454
rect 10208 291134 10528 291218
rect 10208 290898 10250 291134
rect 10486 290898 10528 291134
rect 10208 290866 10528 290898
rect 40928 291454 41248 291486
rect 40928 291218 40970 291454
rect 41206 291218 41248 291454
rect 40928 291134 41248 291218
rect 40928 290898 40970 291134
rect 41206 290898 41248 291134
rect 40928 290866 41248 290898
rect 71648 291454 71968 291486
rect 71648 291218 71690 291454
rect 71926 291218 71968 291454
rect 71648 291134 71968 291218
rect 71648 290898 71690 291134
rect 71926 290898 71968 291134
rect 71648 290866 71968 290898
rect 102368 291454 102688 291486
rect 102368 291218 102410 291454
rect 102646 291218 102688 291454
rect 102368 291134 102688 291218
rect 102368 290898 102410 291134
rect 102646 290898 102688 291134
rect 102368 290866 102688 290898
rect 133088 291454 133408 291486
rect 133088 291218 133130 291454
rect 133366 291218 133408 291454
rect 133088 291134 133408 291218
rect 133088 290898 133130 291134
rect 133366 290898 133408 291134
rect 133088 290866 133408 290898
rect 163808 291454 164128 291486
rect 163808 291218 163850 291454
rect 164086 291218 164128 291454
rect 163808 291134 164128 291218
rect 163808 290898 163850 291134
rect 164086 290898 164128 291134
rect 163808 290866 164128 290898
rect 194528 291454 194848 291486
rect 194528 291218 194570 291454
rect 194806 291218 194848 291454
rect 194528 291134 194848 291218
rect 194528 290898 194570 291134
rect 194806 290898 194848 291134
rect 194528 290866 194848 290898
rect 225248 291454 225568 291486
rect 225248 291218 225290 291454
rect 225526 291218 225568 291454
rect 225248 291134 225568 291218
rect 225248 290898 225290 291134
rect 225526 290898 225568 291134
rect 225248 290866 225568 290898
rect 255968 291454 256288 291486
rect 255968 291218 256010 291454
rect 256246 291218 256288 291454
rect 255968 291134 256288 291218
rect 255968 290898 256010 291134
rect 256246 290898 256288 291134
rect 255968 290866 256288 290898
rect 286688 291454 287008 291486
rect 286688 291218 286730 291454
rect 286966 291218 287008 291454
rect 286688 291134 287008 291218
rect 286688 290898 286730 291134
rect 286966 290898 287008 291134
rect 286688 290866 287008 290898
rect 317408 291454 317728 291486
rect 317408 291218 317450 291454
rect 317686 291218 317728 291454
rect 317408 291134 317728 291218
rect 317408 290898 317450 291134
rect 317686 290898 317728 291134
rect 317408 290866 317728 290898
rect 348128 291454 348448 291486
rect 348128 291218 348170 291454
rect 348406 291218 348448 291454
rect 348128 291134 348448 291218
rect 348128 290898 348170 291134
rect 348406 290898 348448 291134
rect 348128 290866 348448 290898
rect 378848 291454 379168 291486
rect 378848 291218 378890 291454
rect 379126 291218 379168 291454
rect 378848 291134 379168 291218
rect 378848 290898 378890 291134
rect 379126 290898 379168 291134
rect 378848 290866 379168 290898
rect 409568 291454 409888 291486
rect 409568 291218 409610 291454
rect 409846 291218 409888 291454
rect 409568 291134 409888 291218
rect 409568 290898 409610 291134
rect 409846 290898 409888 291134
rect 409568 290866 409888 290898
rect 440288 291454 440608 291486
rect 440288 291218 440330 291454
rect 440566 291218 440608 291454
rect 440288 291134 440608 291218
rect 440288 290898 440330 291134
rect 440566 290898 440608 291134
rect 440288 290866 440608 290898
rect 471008 291454 471328 291486
rect 471008 291218 471050 291454
rect 471286 291218 471328 291454
rect 471008 291134 471328 291218
rect 471008 290898 471050 291134
rect 471286 290898 471328 291134
rect 471008 290866 471328 290898
rect 501728 291454 502048 291486
rect 501728 291218 501770 291454
rect 502006 291218 502048 291454
rect 501728 291134 502048 291218
rect 501728 290898 501770 291134
rect 502006 290898 502048 291134
rect 501728 290866 502048 290898
rect 532448 291454 532768 291486
rect 532448 291218 532490 291454
rect 532726 291218 532768 291454
rect 532448 291134 532768 291218
rect 532448 290898 532490 291134
rect 532726 290898 532768 291134
rect 532448 290866 532768 290898
rect 563168 291454 563488 291486
rect 563168 291218 563210 291454
rect 563446 291218 563488 291454
rect 563168 291134 563488 291218
rect 563168 290898 563210 291134
rect 563446 290898 563488 291134
rect 563168 290866 563488 290898
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 25568 259174 25888 259206
rect 25568 258938 25610 259174
rect 25846 258938 25888 259174
rect 25568 258854 25888 258938
rect 25568 258618 25610 258854
rect 25846 258618 25888 258854
rect 25568 258586 25888 258618
rect 56288 259174 56608 259206
rect 56288 258938 56330 259174
rect 56566 258938 56608 259174
rect 56288 258854 56608 258938
rect 56288 258618 56330 258854
rect 56566 258618 56608 258854
rect 56288 258586 56608 258618
rect 87008 259174 87328 259206
rect 87008 258938 87050 259174
rect 87286 258938 87328 259174
rect 87008 258854 87328 258938
rect 87008 258618 87050 258854
rect 87286 258618 87328 258854
rect 87008 258586 87328 258618
rect 117728 259174 118048 259206
rect 117728 258938 117770 259174
rect 118006 258938 118048 259174
rect 117728 258854 118048 258938
rect 117728 258618 117770 258854
rect 118006 258618 118048 258854
rect 117728 258586 118048 258618
rect 148448 259174 148768 259206
rect 148448 258938 148490 259174
rect 148726 258938 148768 259174
rect 148448 258854 148768 258938
rect 148448 258618 148490 258854
rect 148726 258618 148768 258854
rect 148448 258586 148768 258618
rect 179168 259174 179488 259206
rect 179168 258938 179210 259174
rect 179446 258938 179488 259174
rect 179168 258854 179488 258938
rect 179168 258618 179210 258854
rect 179446 258618 179488 258854
rect 179168 258586 179488 258618
rect 209888 259174 210208 259206
rect 209888 258938 209930 259174
rect 210166 258938 210208 259174
rect 209888 258854 210208 258938
rect 209888 258618 209930 258854
rect 210166 258618 210208 258854
rect 209888 258586 210208 258618
rect 240608 259174 240928 259206
rect 240608 258938 240650 259174
rect 240886 258938 240928 259174
rect 240608 258854 240928 258938
rect 240608 258618 240650 258854
rect 240886 258618 240928 258854
rect 240608 258586 240928 258618
rect 271328 259174 271648 259206
rect 271328 258938 271370 259174
rect 271606 258938 271648 259174
rect 271328 258854 271648 258938
rect 271328 258618 271370 258854
rect 271606 258618 271648 258854
rect 271328 258586 271648 258618
rect 302048 259174 302368 259206
rect 302048 258938 302090 259174
rect 302326 258938 302368 259174
rect 302048 258854 302368 258938
rect 302048 258618 302090 258854
rect 302326 258618 302368 258854
rect 302048 258586 302368 258618
rect 332768 259174 333088 259206
rect 332768 258938 332810 259174
rect 333046 258938 333088 259174
rect 332768 258854 333088 258938
rect 332768 258618 332810 258854
rect 333046 258618 333088 258854
rect 332768 258586 333088 258618
rect 363488 259174 363808 259206
rect 363488 258938 363530 259174
rect 363766 258938 363808 259174
rect 363488 258854 363808 258938
rect 363488 258618 363530 258854
rect 363766 258618 363808 258854
rect 363488 258586 363808 258618
rect 394208 259174 394528 259206
rect 394208 258938 394250 259174
rect 394486 258938 394528 259174
rect 394208 258854 394528 258938
rect 394208 258618 394250 258854
rect 394486 258618 394528 258854
rect 394208 258586 394528 258618
rect 424928 259174 425248 259206
rect 424928 258938 424970 259174
rect 425206 258938 425248 259174
rect 424928 258854 425248 258938
rect 424928 258618 424970 258854
rect 425206 258618 425248 258854
rect 424928 258586 425248 258618
rect 455648 259174 455968 259206
rect 455648 258938 455690 259174
rect 455926 258938 455968 259174
rect 455648 258854 455968 258938
rect 455648 258618 455690 258854
rect 455926 258618 455968 258854
rect 455648 258586 455968 258618
rect 486368 259174 486688 259206
rect 486368 258938 486410 259174
rect 486646 258938 486688 259174
rect 486368 258854 486688 258938
rect 486368 258618 486410 258854
rect 486646 258618 486688 258854
rect 486368 258586 486688 258618
rect 517088 259174 517408 259206
rect 517088 258938 517130 259174
rect 517366 258938 517408 259174
rect 517088 258854 517408 258938
rect 517088 258618 517130 258854
rect 517366 258618 517408 258854
rect 517088 258586 517408 258618
rect 547808 259174 548128 259206
rect 547808 258938 547850 259174
rect 548086 258938 548128 259174
rect 547808 258854 548128 258938
rect 547808 258618 547850 258854
rect 548086 258618 548128 258854
rect 547808 258586 548128 258618
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 10208 255454 10528 255486
rect 10208 255218 10250 255454
rect 10486 255218 10528 255454
rect 10208 255134 10528 255218
rect 10208 254898 10250 255134
rect 10486 254898 10528 255134
rect 10208 254866 10528 254898
rect 40928 255454 41248 255486
rect 40928 255218 40970 255454
rect 41206 255218 41248 255454
rect 40928 255134 41248 255218
rect 40928 254898 40970 255134
rect 41206 254898 41248 255134
rect 40928 254866 41248 254898
rect 71648 255454 71968 255486
rect 71648 255218 71690 255454
rect 71926 255218 71968 255454
rect 71648 255134 71968 255218
rect 71648 254898 71690 255134
rect 71926 254898 71968 255134
rect 71648 254866 71968 254898
rect 102368 255454 102688 255486
rect 102368 255218 102410 255454
rect 102646 255218 102688 255454
rect 102368 255134 102688 255218
rect 102368 254898 102410 255134
rect 102646 254898 102688 255134
rect 102368 254866 102688 254898
rect 133088 255454 133408 255486
rect 133088 255218 133130 255454
rect 133366 255218 133408 255454
rect 133088 255134 133408 255218
rect 133088 254898 133130 255134
rect 133366 254898 133408 255134
rect 133088 254866 133408 254898
rect 163808 255454 164128 255486
rect 163808 255218 163850 255454
rect 164086 255218 164128 255454
rect 163808 255134 164128 255218
rect 163808 254898 163850 255134
rect 164086 254898 164128 255134
rect 163808 254866 164128 254898
rect 194528 255454 194848 255486
rect 194528 255218 194570 255454
rect 194806 255218 194848 255454
rect 194528 255134 194848 255218
rect 194528 254898 194570 255134
rect 194806 254898 194848 255134
rect 194528 254866 194848 254898
rect 225248 255454 225568 255486
rect 225248 255218 225290 255454
rect 225526 255218 225568 255454
rect 225248 255134 225568 255218
rect 225248 254898 225290 255134
rect 225526 254898 225568 255134
rect 225248 254866 225568 254898
rect 255968 255454 256288 255486
rect 255968 255218 256010 255454
rect 256246 255218 256288 255454
rect 255968 255134 256288 255218
rect 255968 254898 256010 255134
rect 256246 254898 256288 255134
rect 255968 254866 256288 254898
rect 286688 255454 287008 255486
rect 286688 255218 286730 255454
rect 286966 255218 287008 255454
rect 286688 255134 287008 255218
rect 286688 254898 286730 255134
rect 286966 254898 287008 255134
rect 286688 254866 287008 254898
rect 317408 255454 317728 255486
rect 317408 255218 317450 255454
rect 317686 255218 317728 255454
rect 317408 255134 317728 255218
rect 317408 254898 317450 255134
rect 317686 254898 317728 255134
rect 317408 254866 317728 254898
rect 348128 255454 348448 255486
rect 348128 255218 348170 255454
rect 348406 255218 348448 255454
rect 348128 255134 348448 255218
rect 348128 254898 348170 255134
rect 348406 254898 348448 255134
rect 348128 254866 348448 254898
rect 378848 255454 379168 255486
rect 378848 255218 378890 255454
rect 379126 255218 379168 255454
rect 378848 255134 379168 255218
rect 378848 254898 378890 255134
rect 379126 254898 379168 255134
rect 378848 254866 379168 254898
rect 409568 255454 409888 255486
rect 409568 255218 409610 255454
rect 409846 255218 409888 255454
rect 409568 255134 409888 255218
rect 409568 254898 409610 255134
rect 409846 254898 409888 255134
rect 409568 254866 409888 254898
rect 440288 255454 440608 255486
rect 440288 255218 440330 255454
rect 440566 255218 440608 255454
rect 440288 255134 440608 255218
rect 440288 254898 440330 255134
rect 440566 254898 440608 255134
rect 440288 254866 440608 254898
rect 471008 255454 471328 255486
rect 471008 255218 471050 255454
rect 471286 255218 471328 255454
rect 471008 255134 471328 255218
rect 471008 254898 471050 255134
rect 471286 254898 471328 255134
rect 471008 254866 471328 254898
rect 501728 255454 502048 255486
rect 501728 255218 501770 255454
rect 502006 255218 502048 255454
rect 501728 255134 502048 255218
rect 501728 254898 501770 255134
rect 502006 254898 502048 255134
rect 501728 254866 502048 254898
rect 532448 255454 532768 255486
rect 532448 255218 532490 255454
rect 532726 255218 532768 255454
rect 532448 255134 532768 255218
rect 532448 254898 532490 255134
rect 532726 254898 532768 255134
rect 532448 254866 532768 254898
rect 563168 255454 563488 255486
rect 563168 255218 563210 255454
rect 563446 255218 563488 255454
rect 563168 255134 563488 255218
rect 563168 254898 563210 255134
rect 563446 254898 563488 255134
rect 563168 254866 563488 254898
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 25568 223174 25888 223206
rect 25568 222938 25610 223174
rect 25846 222938 25888 223174
rect 25568 222854 25888 222938
rect 25568 222618 25610 222854
rect 25846 222618 25888 222854
rect 25568 222586 25888 222618
rect 56288 223174 56608 223206
rect 56288 222938 56330 223174
rect 56566 222938 56608 223174
rect 56288 222854 56608 222938
rect 56288 222618 56330 222854
rect 56566 222618 56608 222854
rect 56288 222586 56608 222618
rect 87008 223174 87328 223206
rect 87008 222938 87050 223174
rect 87286 222938 87328 223174
rect 87008 222854 87328 222938
rect 87008 222618 87050 222854
rect 87286 222618 87328 222854
rect 87008 222586 87328 222618
rect 117728 223174 118048 223206
rect 117728 222938 117770 223174
rect 118006 222938 118048 223174
rect 117728 222854 118048 222938
rect 117728 222618 117770 222854
rect 118006 222618 118048 222854
rect 117728 222586 118048 222618
rect 148448 223174 148768 223206
rect 148448 222938 148490 223174
rect 148726 222938 148768 223174
rect 148448 222854 148768 222938
rect 148448 222618 148490 222854
rect 148726 222618 148768 222854
rect 148448 222586 148768 222618
rect 179168 223174 179488 223206
rect 179168 222938 179210 223174
rect 179446 222938 179488 223174
rect 179168 222854 179488 222938
rect 179168 222618 179210 222854
rect 179446 222618 179488 222854
rect 179168 222586 179488 222618
rect 209888 223174 210208 223206
rect 209888 222938 209930 223174
rect 210166 222938 210208 223174
rect 209888 222854 210208 222938
rect 209888 222618 209930 222854
rect 210166 222618 210208 222854
rect 209888 222586 210208 222618
rect 240608 223174 240928 223206
rect 240608 222938 240650 223174
rect 240886 222938 240928 223174
rect 240608 222854 240928 222938
rect 240608 222618 240650 222854
rect 240886 222618 240928 222854
rect 240608 222586 240928 222618
rect 271328 223174 271648 223206
rect 271328 222938 271370 223174
rect 271606 222938 271648 223174
rect 271328 222854 271648 222938
rect 271328 222618 271370 222854
rect 271606 222618 271648 222854
rect 271328 222586 271648 222618
rect 302048 223174 302368 223206
rect 302048 222938 302090 223174
rect 302326 222938 302368 223174
rect 302048 222854 302368 222938
rect 302048 222618 302090 222854
rect 302326 222618 302368 222854
rect 302048 222586 302368 222618
rect 332768 223174 333088 223206
rect 332768 222938 332810 223174
rect 333046 222938 333088 223174
rect 332768 222854 333088 222938
rect 332768 222618 332810 222854
rect 333046 222618 333088 222854
rect 332768 222586 333088 222618
rect 363488 223174 363808 223206
rect 363488 222938 363530 223174
rect 363766 222938 363808 223174
rect 363488 222854 363808 222938
rect 363488 222618 363530 222854
rect 363766 222618 363808 222854
rect 363488 222586 363808 222618
rect 394208 223174 394528 223206
rect 394208 222938 394250 223174
rect 394486 222938 394528 223174
rect 394208 222854 394528 222938
rect 394208 222618 394250 222854
rect 394486 222618 394528 222854
rect 394208 222586 394528 222618
rect 424928 223174 425248 223206
rect 424928 222938 424970 223174
rect 425206 222938 425248 223174
rect 424928 222854 425248 222938
rect 424928 222618 424970 222854
rect 425206 222618 425248 222854
rect 424928 222586 425248 222618
rect 455648 223174 455968 223206
rect 455648 222938 455690 223174
rect 455926 222938 455968 223174
rect 455648 222854 455968 222938
rect 455648 222618 455690 222854
rect 455926 222618 455968 222854
rect 455648 222586 455968 222618
rect 486368 223174 486688 223206
rect 486368 222938 486410 223174
rect 486646 222938 486688 223174
rect 486368 222854 486688 222938
rect 486368 222618 486410 222854
rect 486646 222618 486688 222854
rect 486368 222586 486688 222618
rect 517088 223174 517408 223206
rect 517088 222938 517130 223174
rect 517366 222938 517408 223174
rect 517088 222854 517408 222938
rect 517088 222618 517130 222854
rect 517366 222618 517408 222854
rect 517088 222586 517408 222618
rect 547808 223174 548128 223206
rect 547808 222938 547850 223174
rect 548086 222938 548128 223174
rect 547808 222854 548128 222938
rect 547808 222618 547850 222854
rect 548086 222618 548128 222854
rect 547808 222586 548128 222618
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 10208 219454 10528 219486
rect 10208 219218 10250 219454
rect 10486 219218 10528 219454
rect 10208 219134 10528 219218
rect 10208 218898 10250 219134
rect 10486 218898 10528 219134
rect 10208 218866 10528 218898
rect 40928 219454 41248 219486
rect 40928 219218 40970 219454
rect 41206 219218 41248 219454
rect 40928 219134 41248 219218
rect 40928 218898 40970 219134
rect 41206 218898 41248 219134
rect 40928 218866 41248 218898
rect 71648 219454 71968 219486
rect 71648 219218 71690 219454
rect 71926 219218 71968 219454
rect 71648 219134 71968 219218
rect 71648 218898 71690 219134
rect 71926 218898 71968 219134
rect 71648 218866 71968 218898
rect 102368 219454 102688 219486
rect 102368 219218 102410 219454
rect 102646 219218 102688 219454
rect 102368 219134 102688 219218
rect 102368 218898 102410 219134
rect 102646 218898 102688 219134
rect 102368 218866 102688 218898
rect 133088 219454 133408 219486
rect 133088 219218 133130 219454
rect 133366 219218 133408 219454
rect 133088 219134 133408 219218
rect 133088 218898 133130 219134
rect 133366 218898 133408 219134
rect 133088 218866 133408 218898
rect 163808 219454 164128 219486
rect 163808 219218 163850 219454
rect 164086 219218 164128 219454
rect 163808 219134 164128 219218
rect 163808 218898 163850 219134
rect 164086 218898 164128 219134
rect 163808 218866 164128 218898
rect 194528 219454 194848 219486
rect 194528 219218 194570 219454
rect 194806 219218 194848 219454
rect 194528 219134 194848 219218
rect 194528 218898 194570 219134
rect 194806 218898 194848 219134
rect 194528 218866 194848 218898
rect 225248 219454 225568 219486
rect 225248 219218 225290 219454
rect 225526 219218 225568 219454
rect 225248 219134 225568 219218
rect 225248 218898 225290 219134
rect 225526 218898 225568 219134
rect 225248 218866 225568 218898
rect 255968 219454 256288 219486
rect 255968 219218 256010 219454
rect 256246 219218 256288 219454
rect 255968 219134 256288 219218
rect 255968 218898 256010 219134
rect 256246 218898 256288 219134
rect 255968 218866 256288 218898
rect 286688 219454 287008 219486
rect 286688 219218 286730 219454
rect 286966 219218 287008 219454
rect 286688 219134 287008 219218
rect 286688 218898 286730 219134
rect 286966 218898 287008 219134
rect 286688 218866 287008 218898
rect 317408 219454 317728 219486
rect 317408 219218 317450 219454
rect 317686 219218 317728 219454
rect 317408 219134 317728 219218
rect 317408 218898 317450 219134
rect 317686 218898 317728 219134
rect 317408 218866 317728 218898
rect 348128 219454 348448 219486
rect 348128 219218 348170 219454
rect 348406 219218 348448 219454
rect 348128 219134 348448 219218
rect 348128 218898 348170 219134
rect 348406 218898 348448 219134
rect 348128 218866 348448 218898
rect 378848 219454 379168 219486
rect 378848 219218 378890 219454
rect 379126 219218 379168 219454
rect 378848 219134 379168 219218
rect 378848 218898 378890 219134
rect 379126 218898 379168 219134
rect 378848 218866 379168 218898
rect 409568 219454 409888 219486
rect 409568 219218 409610 219454
rect 409846 219218 409888 219454
rect 409568 219134 409888 219218
rect 409568 218898 409610 219134
rect 409846 218898 409888 219134
rect 409568 218866 409888 218898
rect 440288 219454 440608 219486
rect 440288 219218 440330 219454
rect 440566 219218 440608 219454
rect 440288 219134 440608 219218
rect 440288 218898 440330 219134
rect 440566 218898 440608 219134
rect 440288 218866 440608 218898
rect 471008 219454 471328 219486
rect 471008 219218 471050 219454
rect 471286 219218 471328 219454
rect 471008 219134 471328 219218
rect 471008 218898 471050 219134
rect 471286 218898 471328 219134
rect 471008 218866 471328 218898
rect 501728 219454 502048 219486
rect 501728 219218 501770 219454
rect 502006 219218 502048 219454
rect 501728 219134 502048 219218
rect 501728 218898 501770 219134
rect 502006 218898 502048 219134
rect 501728 218866 502048 218898
rect 532448 219454 532768 219486
rect 532448 219218 532490 219454
rect 532726 219218 532768 219454
rect 532448 219134 532768 219218
rect 532448 218898 532490 219134
rect 532726 218898 532768 219134
rect 532448 218866 532768 218898
rect 563168 219454 563488 219486
rect 563168 219218 563210 219454
rect 563446 219218 563488 219454
rect 563168 219134 563488 219218
rect 563168 218898 563210 219134
rect 563446 218898 563488 219134
rect 563168 218866 563488 218898
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 25568 187174 25888 187206
rect 25568 186938 25610 187174
rect 25846 186938 25888 187174
rect 25568 186854 25888 186938
rect 25568 186618 25610 186854
rect 25846 186618 25888 186854
rect 25568 186586 25888 186618
rect 56288 187174 56608 187206
rect 56288 186938 56330 187174
rect 56566 186938 56608 187174
rect 56288 186854 56608 186938
rect 56288 186618 56330 186854
rect 56566 186618 56608 186854
rect 56288 186586 56608 186618
rect 87008 187174 87328 187206
rect 87008 186938 87050 187174
rect 87286 186938 87328 187174
rect 87008 186854 87328 186938
rect 87008 186618 87050 186854
rect 87286 186618 87328 186854
rect 87008 186586 87328 186618
rect 117728 187174 118048 187206
rect 117728 186938 117770 187174
rect 118006 186938 118048 187174
rect 117728 186854 118048 186938
rect 117728 186618 117770 186854
rect 118006 186618 118048 186854
rect 117728 186586 118048 186618
rect 148448 187174 148768 187206
rect 148448 186938 148490 187174
rect 148726 186938 148768 187174
rect 148448 186854 148768 186938
rect 148448 186618 148490 186854
rect 148726 186618 148768 186854
rect 148448 186586 148768 186618
rect 179168 187174 179488 187206
rect 179168 186938 179210 187174
rect 179446 186938 179488 187174
rect 179168 186854 179488 186938
rect 179168 186618 179210 186854
rect 179446 186618 179488 186854
rect 179168 186586 179488 186618
rect 209888 187174 210208 187206
rect 209888 186938 209930 187174
rect 210166 186938 210208 187174
rect 209888 186854 210208 186938
rect 209888 186618 209930 186854
rect 210166 186618 210208 186854
rect 209888 186586 210208 186618
rect 240608 187174 240928 187206
rect 240608 186938 240650 187174
rect 240886 186938 240928 187174
rect 240608 186854 240928 186938
rect 240608 186618 240650 186854
rect 240886 186618 240928 186854
rect 240608 186586 240928 186618
rect 271328 187174 271648 187206
rect 271328 186938 271370 187174
rect 271606 186938 271648 187174
rect 271328 186854 271648 186938
rect 271328 186618 271370 186854
rect 271606 186618 271648 186854
rect 271328 186586 271648 186618
rect 302048 187174 302368 187206
rect 302048 186938 302090 187174
rect 302326 186938 302368 187174
rect 302048 186854 302368 186938
rect 302048 186618 302090 186854
rect 302326 186618 302368 186854
rect 302048 186586 302368 186618
rect 332768 187174 333088 187206
rect 332768 186938 332810 187174
rect 333046 186938 333088 187174
rect 332768 186854 333088 186938
rect 332768 186618 332810 186854
rect 333046 186618 333088 186854
rect 332768 186586 333088 186618
rect 363488 187174 363808 187206
rect 363488 186938 363530 187174
rect 363766 186938 363808 187174
rect 363488 186854 363808 186938
rect 363488 186618 363530 186854
rect 363766 186618 363808 186854
rect 363488 186586 363808 186618
rect 394208 187174 394528 187206
rect 394208 186938 394250 187174
rect 394486 186938 394528 187174
rect 394208 186854 394528 186938
rect 394208 186618 394250 186854
rect 394486 186618 394528 186854
rect 394208 186586 394528 186618
rect 424928 187174 425248 187206
rect 424928 186938 424970 187174
rect 425206 186938 425248 187174
rect 424928 186854 425248 186938
rect 424928 186618 424970 186854
rect 425206 186618 425248 186854
rect 424928 186586 425248 186618
rect 455648 187174 455968 187206
rect 455648 186938 455690 187174
rect 455926 186938 455968 187174
rect 455648 186854 455968 186938
rect 455648 186618 455690 186854
rect 455926 186618 455968 186854
rect 455648 186586 455968 186618
rect 486368 187174 486688 187206
rect 486368 186938 486410 187174
rect 486646 186938 486688 187174
rect 486368 186854 486688 186938
rect 486368 186618 486410 186854
rect 486646 186618 486688 186854
rect 486368 186586 486688 186618
rect 517088 187174 517408 187206
rect 517088 186938 517130 187174
rect 517366 186938 517408 187174
rect 517088 186854 517408 186938
rect 517088 186618 517130 186854
rect 517366 186618 517408 186854
rect 517088 186586 517408 186618
rect 547808 187174 548128 187206
rect 547808 186938 547850 187174
rect 548086 186938 548128 187174
rect 547808 186854 548128 186938
rect 547808 186618 547850 186854
rect 548086 186618 548128 186854
rect 547808 186586 548128 186618
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 10208 183454 10528 183486
rect 10208 183218 10250 183454
rect 10486 183218 10528 183454
rect 10208 183134 10528 183218
rect 10208 182898 10250 183134
rect 10486 182898 10528 183134
rect 10208 182866 10528 182898
rect 40928 183454 41248 183486
rect 40928 183218 40970 183454
rect 41206 183218 41248 183454
rect 40928 183134 41248 183218
rect 40928 182898 40970 183134
rect 41206 182898 41248 183134
rect 40928 182866 41248 182898
rect 71648 183454 71968 183486
rect 71648 183218 71690 183454
rect 71926 183218 71968 183454
rect 71648 183134 71968 183218
rect 71648 182898 71690 183134
rect 71926 182898 71968 183134
rect 71648 182866 71968 182898
rect 102368 183454 102688 183486
rect 102368 183218 102410 183454
rect 102646 183218 102688 183454
rect 102368 183134 102688 183218
rect 102368 182898 102410 183134
rect 102646 182898 102688 183134
rect 102368 182866 102688 182898
rect 133088 183454 133408 183486
rect 133088 183218 133130 183454
rect 133366 183218 133408 183454
rect 133088 183134 133408 183218
rect 133088 182898 133130 183134
rect 133366 182898 133408 183134
rect 133088 182866 133408 182898
rect 163808 183454 164128 183486
rect 163808 183218 163850 183454
rect 164086 183218 164128 183454
rect 163808 183134 164128 183218
rect 163808 182898 163850 183134
rect 164086 182898 164128 183134
rect 163808 182866 164128 182898
rect 194528 183454 194848 183486
rect 194528 183218 194570 183454
rect 194806 183218 194848 183454
rect 194528 183134 194848 183218
rect 194528 182898 194570 183134
rect 194806 182898 194848 183134
rect 194528 182866 194848 182898
rect 225248 183454 225568 183486
rect 225248 183218 225290 183454
rect 225526 183218 225568 183454
rect 225248 183134 225568 183218
rect 225248 182898 225290 183134
rect 225526 182898 225568 183134
rect 225248 182866 225568 182898
rect 255968 183454 256288 183486
rect 255968 183218 256010 183454
rect 256246 183218 256288 183454
rect 255968 183134 256288 183218
rect 255968 182898 256010 183134
rect 256246 182898 256288 183134
rect 255968 182866 256288 182898
rect 286688 183454 287008 183486
rect 286688 183218 286730 183454
rect 286966 183218 287008 183454
rect 286688 183134 287008 183218
rect 286688 182898 286730 183134
rect 286966 182898 287008 183134
rect 286688 182866 287008 182898
rect 317408 183454 317728 183486
rect 317408 183218 317450 183454
rect 317686 183218 317728 183454
rect 317408 183134 317728 183218
rect 317408 182898 317450 183134
rect 317686 182898 317728 183134
rect 317408 182866 317728 182898
rect 348128 183454 348448 183486
rect 348128 183218 348170 183454
rect 348406 183218 348448 183454
rect 348128 183134 348448 183218
rect 348128 182898 348170 183134
rect 348406 182898 348448 183134
rect 348128 182866 348448 182898
rect 378848 183454 379168 183486
rect 378848 183218 378890 183454
rect 379126 183218 379168 183454
rect 378848 183134 379168 183218
rect 378848 182898 378890 183134
rect 379126 182898 379168 183134
rect 378848 182866 379168 182898
rect 409568 183454 409888 183486
rect 409568 183218 409610 183454
rect 409846 183218 409888 183454
rect 409568 183134 409888 183218
rect 409568 182898 409610 183134
rect 409846 182898 409888 183134
rect 409568 182866 409888 182898
rect 440288 183454 440608 183486
rect 440288 183218 440330 183454
rect 440566 183218 440608 183454
rect 440288 183134 440608 183218
rect 440288 182898 440330 183134
rect 440566 182898 440608 183134
rect 440288 182866 440608 182898
rect 471008 183454 471328 183486
rect 471008 183218 471050 183454
rect 471286 183218 471328 183454
rect 471008 183134 471328 183218
rect 471008 182898 471050 183134
rect 471286 182898 471328 183134
rect 471008 182866 471328 182898
rect 501728 183454 502048 183486
rect 501728 183218 501770 183454
rect 502006 183218 502048 183454
rect 501728 183134 502048 183218
rect 501728 182898 501770 183134
rect 502006 182898 502048 183134
rect 501728 182866 502048 182898
rect 532448 183454 532768 183486
rect 532448 183218 532490 183454
rect 532726 183218 532768 183454
rect 532448 183134 532768 183218
rect 532448 182898 532490 183134
rect 532726 182898 532768 183134
rect 532448 182866 532768 182898
rect 563168 183454 563488 183486
rect 563168 183218 563210 183454
rect 563446 183218 563488 183454
rect 563168 183134 563488 183218
rect 563168 182898 563210 183134
rect 563446 182898 563488 183134
rect 563168 182866 563488 182898
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 25568 151174 25888 151206
rect 25568 150938 25610 151174
rect 25846 150938 25888 151174
rect 25568 150854 25888 150938
rect 25568 150618 25610 150854
rect 25846 150618 25888 150854
rect 25568 150586 25888 150618
rect 56288 151174 56608 151206
rect 56288 150938 56330 151174
rect 56566 150938 56608 151174
rect 56288 150854 56608 150938
rect 56288 150618 56330 150854
rect 56566 150618 56608 150854
rect 56288 150586 56608 150618
rect 87008 151174 87328 151206
rect 87008 150938 87050 151174
rect 87286 150938 87328 151174
rect 87008 150854 87328 150938
rect 87008 150618 87050 150854
rect 87286 150618 87328 150854
rect 87008 150586 87328 150618
rect 117728 151174 118048 151206
rect 117728 150938 117770 151174
rect 118006 150938 118048 151174
rect 117728 150854 118048 150938
rect 117728 150618 117770 150854
rect 118006 150618 118048 150854
rect 117728 150586 118048 150618
rect 148448 151174 148768 151206
rect 148448 150938 148490 151174
rect 148726 150938 148768 151174
rect 148448 150854 148768 150938
rect 148448 150618 148490 150854
rect 148726 150618 148768 150854
rect 148448 150586 148768 150618
rect 179168 151174 179488 151206
rect 179168 150938 179210 151174
rect 179446 150938 179488 151174
rect 179168 150854 179488 150938
rect 179168 150618 179210 150854
rect 179446 150618 179488 150854
rect 179168 150586 179488 150618
rect 209888 151174 210208 151206
rect 209888 150938 209930 151174
rect 210166 150938 210208 151174
rect 209888 150854 210208 150938
rect 209888 150618 209930 150854
rect 210166 150618 210208 150854
rect 209888 150586 210208 150618
rect 240608 151174 240928 151206
rect 240608 150938 240650 151174
rect 240886 150938 240928 151174
rect 240608 150854 240928 150938
rect 240608 150618 240650 150854
rect 240886 150618 240928 150854
rect 240608 150586 240928 150618
rect 271328 151174 271648 151206
rect 271328 150938 271370 151174
rect 271606 150938 271648 151174
rect 271328 150854 271648 150938
rect 271328 150618 271370 150854
rect 271606 150618 271648 150854
rect 271328 150586 271648 150618
rect 302048 151174 302368 151206
rect 302048 150938 302090 151174
rect 302326 150938 302368 151174
rect 302048 150854 302368 150938
rect 302048 150618 302090 150854
rect 302326 150618 302368 150854
rect 302048 150586 302368 150618
rect 332768 151174 333088 151206
rect 332768 150938 332810 151174
rect 333046 150938 333088 151174
rect 332768 150854 333088 150938
rect 332768 150618 332810 150854
rect 333046 150618 333088 150854
rect 332768 150586 333088 150618
rect 363488 151174 363808 151206
rect 363488 150938 363530 151174
rect 363766 150938 363808 151174
rect 363488 150854 363808 150938
rect 363488 150618 363530 150854
rect 363766 150618 363808 150854
rect 363488 150586 363808 150618
rect 394208 151174 394528 151206
rect 394208 150938 394250 151174
rect 394486 150938 394528 151174
rect 394208 150854 394528 150938
rect 394208 150618 394250 150854
rect 394486 150618 394528 150854
rect 394208 150586 394528 150618
rect 424928 151174 425248 151206
rect 424928 150938 424970 151174
rect 425206 150938 425248 151174
rect 424928 150854 425248 150938
rect 424928 150618 424970 150854
rect 425206 150618 425248 150854
rect 424928 150586 425248 150618
rect 455648 151174 455968 151206
rect 455648 150938 455690 151174
rect 455926 150938 455968 151174
rect 455648 150854 455968 150938
rect 455648 150618 455690 150854
rect 455926 150618 455968 150854
rect 455648 150586 455968 150618
rect 486368 151174 486688 151206
rect 486368 150938 486410 151174
rect 486646 150938 486688 151174
rect 486368 150854 486688 150938
rect 486368 150618 486410 150854
rect 486646 150618 486688 150854
rect 486368 150586 486688 150618
rect 517088 151174 517408 151206
rect 517088 150938 517130 151174
rect 517366 150938 517408 151174
rect 517088 150854 517408 150938
rect 517088 150618 517130 150854
rect 517366 150618 517408 150854
rect 517088 150586 517408 150618
rect 547808 151174 548128 151206
rect 547808 150938 547850 151174
rect 548086 150938 548128 151174
rect 547808 150854 548128 150938
rect 547808 150618 547850 150854
rect 548086 150618 548128 150854
rect 547808 150586 548128 150618
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 10208 147454 10528 147486
rect 10208 147218 10250 147454
rect 10486 147218 10528 147454
rect 10208 147134 10528 147218
rect 10208 146898 10250 147134
rect 10486 146898 10528 147134
rect 10208 146866 10528 146898
rect 40928 147454 41248 147486
rect 40928 147218 40970 147454
rect 41206 147218 41248 147454
rect 40928 147134 41248 147218
rect 40928 146898 40970 147134
rect 41206 146898 41248 147134
rect 40928 146866 41248 146898
rect 71648 147454 71968 147486
rect 71648 147218 71690 147454
rect 71926 147218 71968 147454
rect 71648 147134 71968 147218
rect 71648 146898 71690 147134
rect 71926 146898 71968 147134
rect 71648 146866 71968 146898
rect 102368 147454 102688 147486
rect 102368 147218 102410 147454
rect 102646 147218 102688 147454
rect 102368 147134 102688 147218
rect 102368 146898 102410 147134
rect 102646 146898 102688 147134
rect 102368 146866 102688 146898
rect 133088 147454 133408 147486
rect 133088 147218 133130 147454
rect 133366 147218 133408 147454
rect 133088 147134 133408 147218
rect 133088 146898 133130 147134
rect 133366 146898 133408 147134
rect 133088 146866 133408 146898
rect 163808 147454 164128 147486
rect 163808 147218 163850 147454
rect 164086 147218 164128 147454
rect 163808 147134 164128 147218
rect 163808 146898 163850 147134
rect 164086 146898 164128 147134
rect 163808 146866 164128 146898
rect 194528 147454 194848 147486
rect 194528 147218 194570 147454
rect 194806 147218 194848 147454
rect 194528 147134 194848 147218
rect 194528 146898 194570 147134
rect 194806 146898 194848 147134
rect 194528 146866 194848 146898
rect 225248 147454 225568 147486
rect 225248 147218 225290 147454
rect 225526 147218 225568 147454
rect 225248 147134 225568 147218
rect 225248 146898 225290 147134
rect 225526 146898 225568 147134
rect 225248 146866 225568 146898
rect 255968 147454 256288 147486
rect 255968 147218 256010 147454
rect 256246 147218 256288 147454
rect 255968 147134 256288 147218
rect 255968 146898 256010 147134
rect 256246 146898 256288 147134
rect 255968 146866 256288 146898
rect 286688 147454 287008 147486
rect 286688 147218 286730 147454
rect 286966 147218 287008 147454
rect 286688 147134 287008 147218
rect 286688 146898 286730 147134
rect 286966 146898 287008 147134
rect 286688 146866 287008 146898
rect 317408 147454 317728 147486
rect 317408 147218 317450 147454
rect 317686 147218 317728 147454
rect 317408 147134 317728 147218
rect 317408 146898 317450 147134
rect 317686 146898 317728 147134
rect 317408 146866 317728 146898
rect 348128 147454 348448 147486
rect 348128 147218 348170 147454
rect 348406 147218 348448 147454
rect 348128 147134 348448 147218
rect 348128 146898 348170 147134
rect 348406 146898 348448 147134
rect 348128 146866 348448 146898
rect 378848 147454 379168 147486
rect 378848 147218 378890 147454
rect 379126 147218 379168 147454
rect 378848 147134 379168 147218
rect 378848 146898 378890 147134
rect 379126 146898 379168 147134
rect 378848 146866 379168 146898
rect 409568 147454 409888 147486
rect 409568 147218 409610 147454
rect 409846 147218 409888 147454
rect 409568 147134 409888 147218
rect 409568 146898 409610 147134
rect 409846 146898 409888 147134
rect 409568 146866 409888 146898
rect 440288 147454 440608 147486
rect 440288 147218 440330 147454
rect 440566 147218 440608 147454
rect 440288 147134 440608 147218
rect 440288 146898 440330 147134
rect 440566 146898 440608 147134
rect 440288 146866 440608 146898
rect 471008 147454 471328 147486
rect 471008 147218 471050 147454
rect 471286 147218 471328 147454
rect 471008 147134 471328 147218
rect 471008 146898 471050 147134
rect 471286 146898 471328 147134
rect 471008 146866 471328 146898
rect 501728 147454 502048 147486
rect 501728 147218 501770 147454
rect 502006 147218 502048 147454
rect 501728 147134 502048 147218
rect 501728 146898 501770 147134
rect 502006 146898 502048 147134
rect 501728 146866 502048 146898
rect 532448 147454 532768 147486
rect 532448 147218 532490 147454
rect 532726 147218 532768 147454
rect 532448 147134 532768 147218
rect 532448 146898 532490 147134
rect 532726 146898 532768 147134
rect 532448 146866 532768 146898
rect 563168 147454 563488 147486
rect 563168 147218 563210 147454
rect 563446 147218 563488 147454
rect 563168 147134 563488 147218
rect 563168 146898 563210 147134
rect 563446 146898 563488 147134
rect 563168 146866 563488 146898
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 25568 115174 25888 115206
rect 25568 114938 25610 115174
rect 25846 114938 25888 115174
rect 25568 114854 25888 114938
rect 25568 114618 25610 114854
rect 25846 114618 25888 114854
rect 25568 114586 25888 114618
rect 56288 115174 56608 115206
rect 56288 114938 56330 115174
rect 56566 114938 56608 115174
rect 56288 114854 56608 114938
rect 56288 114618 56330 114854
rect 56566 114618 56608 114854
rect 56288 114586 56608 114618
rect 87008 115174 87328 115206
rect 87008 114938 87050 115174
rect 87286 114938 87328 115174
rect 87008 114854 87328 114938
rect 87008 114618 87050 114854
rect 87286 114618 87328 114854
rect 87008 114586 87328 114618
rect 117728 115174 118048 115206
rect 117728 114938 117770 115174
rect 118006 114938 118048 115174
rect 117728 114854 118048 114938
rect 117728 114618 117770 114854
rect 118006 114618 118048 114854
rect 117728 114586 118048 114618
rect 148448 115174 148768 115206
rect 148448 114938 148490 115174
rect 148726 114938 148768 115174
rect 148448 114854 148768 114938
rect 148448 114618 148490 114854
rect 148726 114618 148768 114854
rect 148448 114586 148768 114618
rect 179168 115174 179488 115206
rect 179168 114938 179210 115174
rect 179446 114938 179488 115174
rect 179168 114854 179488 114938
rect 179168 114618 179210 114854
rect 179446 114618 179488 114854
rect 179168 114586 179488 114618
rect 209888 115174 210208 115206
rect 209888 114938 209930 115174
rect 210166 114938 210208 115174
rect 209888 114854 210208 114938
rect 209888 114618 209930 114854
rect 210166 114618 210208 114854
rect 209888 114586 210208 114618
rect 240608 115174 240928 115206
rect 240608 114938 240650 115174
rect 240886 114938 240928 115174
rect 240608 114854 240928 114938
rect 240608 114618 240650 114854
rect 240886 114618 240928 114854
rect 240608 114586 240928 114618
rect 271328 115174 271648 115206
rect 271328 114938 271370 115174
rect 271606 114938 271648 115174
rect 271328 114854 271648 114938
rect 271328 114618 271370 114854
rect 271606 114618 271648 114854
rect 271328 114586 271648 114618
rect 302048 115174 302368 115206
rect 302048 114938 302090 115174
rect 302326 114938 302368 115174
rect 302048 114854 302368 114938
rect 302048 114618 302090 114854
rect 302326 114618 302368 114854
rect 302048 114586 302368 114618
rect 332768 115174 333088 115206
rect 332768 114938 332810 115174
rect 333046 114938 333088 115174
rect 332768 114854 333088 114938
rect 332768 114618 332810 114854
rect 333046 114618 333088 114854
rect 332768 114586 333088 114618
rect 363488 115174 363808 115206
rect 363488 114938 363530 115174
rect 363766 114938 363808 115174
rect 363488 114854 363808 114938
rect 363488 114618 363530 114854
rect 363766 114618 363808 114854
rect 363488 114586 363808 114618
rect 394208 115174 394528 115206
rect 394208 114938 394250 115174
rect 394486 114938 394528 115174
rect 394208 114854 394528 114938
rect 394208 114618 394250 114854
rect 394486 114618 394528 114854
rect 394208 114586 394528 114618
rect 424928 115174 425248 115206
rect 424928 114938 424970 115174
rect 425206 114938 425248 115174
rect 424928 114854 425248 114938
rect 424928 114618 424970 114854
rect 425206 114618 425248 114854
rect 424928 114586 425248 114618
rect 455648 115174 455968 115206
rect 455648 114938 455690 115174
rect 455926 114938 455968 115174
rect 455648 114854 455968 114938
rect 455648 114618 455690 114854
rect 455926 114618 455968 114854
rect 455648 114586 455968 114618
rect 486368 115174 486688 115206
rect 486368 114938 486410 115174
rect 486646 114938 486688 115174
rect 486368 114854 486688 114938
rect 486368 114618 486410 114854
rect 486646 114618 486688 114854
rect 486368 114586 486688 114618
rect 517088 115174 517408 115206
rect 517088 114938 517130 115174
rect 517366 114938 517408 115174
rect 517088 114854 517408 114938
rect 517088 114618 517130 114854
rect 517366 114618 517408 114854
rect 517088 114586 517408 114618
rect 547808 115174 548128 115206
rect 547808 114938 547850 115174
rect 548086 114938 548128 115174
rect 547808 114854 548128 114938
rect 547808 114618 547850 114854
rect 548086 114618 548128 114854
rect 547808 114586 548128 114618
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 10208 111454 10528 111486
rect 10208 111218 10250 111454
rect 10486 111218 10528 111454
rect 10208 111134 10528 111218
rect 10208 110898 10250 111134
rect 10486 110898 10528 111134
rect 10208 110866 10528 110898
rect 40928 111454 41248 111486
rect 40928 111218 40970 111454
rect 41206 111218 41248 111454
rect 40928 111134 41248 111218
rect 40928 110898 40970 111134
rect 41206 110898 41248 111134
rect 40928 110866 41248 110898
rect 71648 111454 71968 111486
rect 71648 111218 71690 111454
rect 71926 111218 71968 111454
rect 71648 111134 71968 111218
rect 71648 110898 71690 111134
rect 71926 110898 71968 111134
rect 71648 110866 71968 110898
rect 102368 111454 102688 111486
rect 102368 111218 102410 111454
rect 102646 111218 102688 111454
rect 102368 111134 102688 111218
rect 102368 110898 102410 111134
rect 102646 110898 102688 111134
rect 102368 110866 102688 110898
rect 133088 111454 133408 111486
rect 133088 111218 133130 111454
rect 133366 111218 133408 111454
rect 133088 111134 133408 111218
rect 133088 110898 133130 111134
rect 133366 110898 133408 111134
rect 133088 110866 133408 110898
rect 163808 111454 164128 111486
rect 163808 111218 163850 111454
rect 164086 111218 164128 111454
rect 163808 111134 164128 111218
rect 163808 110898 163850 111134
rect 164086 110898 164128 111134
rect 163808 110866 164128 110898
rect 194528 111454 194848 111486
rect 194528 111218 194570 111454
rect 194806 111218 194848 111454
rect 194528 111134 194848 111218
rect 194528 110898 194570 111134
rect 194806 110898 194848 111134
rect 194528 110866 194848 110898
rect 225248 111454 225568 111486
rect 225248 111218 225290 111454
rect 225526 111218 225568 111454
rect 225248 111134 225568 111218
rect 225248 110898 225290 111134
rect 225526 110898 225568 111134
rect 225248 110866 225568 110898
rect 255968 111454 256288 111486
rect 255968 111218 256010 111454
rect 256246 111218 256288 111454
rect 255968 111134 256288 111218
rect 255968 110898 256010 111134
rect 256246 110898 256288 111134
rect 255968 110866 256288 110898
rect 286688 111454 287008 111486
rect 286688 111218 286730 111454
rect 286966 111218 287008 111454
rect 286688 111134 287008 111218
rect 286688 110898 286730 111134
rect 286966 110898 287008 111134
rect 286688 110866 287008 110898
rect 317408 111454 317728 111486
rect 317408 111218 317450 111454
rect 317686 111218 317728 111454
rect 317408 111134 317728 111218
rect 317408 110898 317450 111134
rect 317686 110898 317728 111134
rect 317408 110866 317728 110898
rect 348128 111454 348448 111486
rect 348128 111218 348170 111454
rect 348406 111218 348448 111454
rect 348128 111134 348448 111218
rect 348128 110898 348170 111134
rect 348406 110898 348448 111134
rect 348128 110866 348448 110898
rect 378848 111454 379168 111486
rect 378848 111218 378890 111454
rect 379126 111218 379168 111454
rect 378848 111134 379168 111218
rect 378848 110898 378890 111134
rect 379126 110898 379168 111134
rect 378848 110866 379168 110898
rect 409568 111454 409888 111486
rect 409568 111218 409610 111454
rect 409846 111218 409888 111454
rect 409568 111134 409888 111218
rect 409568 110898 409610 111134
rect 409846 110898 409888 111134
rect 409568 110866 409888 110898
rect 440288 111454 440608 111486
rect 440288 111218 440330 111454
rect 440566 111218 440608 111454
rect 440288 111134 440608 111218
rect 440288 110898 440330 111134
rect 440566 110898 440608 111134
rect 440288 110866 440608 110898
rect 471008 111454 471328 111486
rect 471008 111218 471050 111454
rect 471286 111218 471328 111454
rect 471008 111134 471328 111218
rect 471008 110898 471050 111134
rect 471286 110898 471328 111134
rect 471008 110866 471328 110898
rect 501728 111454 502048 111486
rect 501728 111218 501770 111454
rect 502006 111218 502048 111454
rect 501728 111134 502048 111218
rect 501728 110898 501770 111134
rect 502006 110898 502048 111134
rect 501728 110866 502048 110898
rect 532448 111454 532768 111486
rect 532448 111218 532490 111454
rect 532726 111218 532768 111454
rect 532448 111134 532768 111218
rect 532448 110898 532490 111134
rect 532726 110898 532768 111134
rect 532448 110866 532768 110898
rect 563168 111454 563488 111486
rect 563168 111218 563210 111454
rect 563446 111218 563488 111454
rect 563168 111134 563488 111218
rect 563168 110898 563210 111134
rect 563446 110898 563488 111134
rect 563168 110866 563488 110898
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 25568 79174 25888 79206
rect 25568 78938 25610 79174
rect 25846 78938 25888 79174
rect 25568 78854 25888 78938
rect 25568 78618 25610 78854
rect 25846 78618 25888 78854
rect 25568 78586 25888 78618
rect 56288 79174 56608 79206
rect 56288 78938 56330 79174
rect 56566 78938 56608 79174
rect 56288 78854 56608 78938
rect 56288 78618 56330 78854
rect 56566 78618 56608 78854
rect 56288 78586 56608 78618
rect 87008 79174 87328 79206
rect 87008 78938 87050 79174
rect 87286 78938 87328 79174
rect 87008 78854 87328 78938
rect 87008 78618 87050 78854
rect 87286 78618 87328 78854
rect 87008 78586 87328 78618
rect 117728 79174 118048 79206
rect 117728 78938 117770 79174
rect 118006 78938 118048 79174
rect 117728 78854 118048 78938
rect 117728 78618 117770 78854
rect 118006 78618 118048 78854
rect 117728 78586 118048 78618
rect 148448 79174 148768 79206
rect 148448 78938 148490 79174
rect 148726 78938 148768 79174
rect 148448 78854 148768 78938
rect 148448 78618 148490 78854
rect 148726 78618 148768 78854
rect 148448 78586 148768 78618
rect 179168 79174 179488 79206
rect 179168 78938 179210 79174
rect 179446 78938 179488 79174
rect 179168 78854 179488 78938
rect 179168 78618 179210 78854
rect 179446 78618 179488 78854
rect 179168 78586 179488 78618
rect 209888 79174 210208 79206
rect 209888 78938 209930 79174
rect 210166 78938 210208 79174
rect 209888 78854 210208 78938
rect 209888 78618 209930 78854
rect 210166 78618 210208 78854
rect 209888 78586 210208 78618
rect 240608 79174 240928 79206
rect 240608 78938 240650 79174
rect 240886 78938 240928 79174
rect 240608 78854 240928 78938
rect 240608 78618 240650 78854
rect 240886 78618 240928 78854
rect 240608 78586 240928 78618
rect 271328 79174 271648 79206
rect 271328 78938 271370 79174
rect 271606 78938 271648 79174
rect 271328 78854 271648 78938
rect 271328 78618 271370 78854
rect 271606 78618 271648 78854
rect 271328 78586 271648 78618
rect 302048 79174 302368 79206
rect 302048 78938 302090 79174
rect 302326 78938 302368 79174
rect 302048 78854 302368 78938
rect 302048 78618 302090 78854
rect 302326 78618 302368 78854
rect 302048 78586 302368 78618
rect 332768 79174 333088 79206
rect 332768 78938 332810 79174
rect 333046 78938 333088 79174
rect 332768 78854 333088 78938
rect 332768 78618 332810 78854
rect 333046 78618 333088 78854
rect 332768 78586 333088 78618
rect 363488 79174 363808 79206
rect 363488 78938 363530 79174
rect 363766 78938 363808 79174
rect 363488 78854 363808 78938
rect 363488 78618 363530 78854
rect 363766 78618 363808 78854
rect 363488 78586 363808 78618
rect 394208 79174 394528 79206
rect 394208 78938 394250 79174
rect 394486 78938 394528 79174
rect 394208 78854 394528 78938
rect 394208 78618 394250 78854
rect 394486 78618 394528 78854
rect 394208 78586 394528 78618
rect 424928 79174 425248 79206
rect 424928 78938 424970 79174
rect 425206 78938 425248 79174
rect 424928 78854 425248 78938
rect 424928 78618 424970 78854
rect 425206 78618 425248 78854
rect 424928 78586 425248 78618
rect 455648 79174 455968 79206
rect 455648 78938 455690 79174
rect 455926 78938 455968 79174
rect 455648 78854 455968 78938
rect 455648 78618 455690 78854
rect 455926 78618 455968 78854
rect 455648 78586 455968 78618
rect 486368 79174 486688 79206
rect 486368 78938 486410 79174
rect 486646 78938 486688 79174
rect 486368 78854 486688 78938
rect 486368 78618 486410 78854
rect 486646 78618 486688 78854
rect 486368 78586 486688 78618
rect 517088 79174 517408 79206
rect 517088 78938 517130 79174
rect 517366 78938 517408 79174
rect 517088 78854 517408 78938
rect 517088 78618 517130 78854
rect 517366 78618 517408 78854
rect 517088 78586 517408 78618
rect 547808 79174 548128 79206
rect 547808 78938 547850 79174
rect 548086 78938 548128 79174
rect 547808 78854 548128 78938
rect 547808 78618 547850 78854
rect 548086 78618 548128 78854
rect 547808 78586 548128 78618
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 10208 75454 10528 75486
rect 10208 75218 10250 75454
rect 10486 75218 10528 75454
rect 10208 75134 10528 75218
rect 10208 74898 10250 75134
rect 10486 74898 10528 75134
rect 10208 74866 10528 74898
rect 40928 75454 41248 75486
rect 40928 75218 40970 75454
rect 41206 75218 41248 75454
rect 40928 75134 41248 75218
rect 40928 74898 40970 75134
rect 41206 74898 41248 75134
rect 40928 74866 41248 74898
rect 71648 75454 71968 75486
rect 71648 75218 71690 75454
rect 71926 75218 71968 75454
rect 71648 75134 71968 75218
rect 71648 74898 71690 75134
rect 71926 74898 71968 75134
rect 71648 74866 71968 74898
rect 102368 75454 102688 75486
rect 102368 75218 102410 75454
rect 102646 75218 102688 75454
rect 102368 75134 102688 75218
rect 102368 74898 102410 75134
rect 102646 74898 102688 75134
rect 102368 74866 102688 74898
rect 133088 75454 133408 75486
rect 133088 75218 133130 75454
rect 133366 75218 133408 75454
rect 133088 75134 133408 75218
rect 133088 74898 133130 75134
rect 133366 74898 133408 75134
rect 133088 74866 133408 74898
rect 163808 75454 164128 75486
rect 163808 75218 163850 75454
rect 164086 75218 164128 75454
rect 163808 75134 164128 75218
rect 163808 74898 163850 75134
rect 164086 74898 164128 75134
rect 163808 74866 164128 74898
rect 194528 75454 194848 75486
rect 194528 75218 194570 75454
rect 194806 75218 194848 75454
rect 194528 75134 194848 75218
rect 194528 74898 194570 75134
rect 194806 74898 194848 75134
rect 194528 74866 194848 74898
rect 225248 75454 225568 75486
rect 225248 75218 225290 75454
rect 225526 75218 225568 75454
rect 225248 75134 225568 75218
rect 225248 74898 225290 75134
rect 225526 74898 225568 75134
rect 225248 74866 225568 74898
rect 255968 75454 256288 75486
rect 255968 75218 256010 75454
rect 256246 75218 256288 75454
rect 255968 75134 256288 75218
rect 255968 74898 256010 75134
rect 256246 74898 256288 75134
rect 255968 74866 256288 74898
rect 286688 75454 287008 75486
rect 286688 75218 286730 75454
rect 286966 75218 287008 75454
rect 286688 75134 287008 75218
rect 286688 74898 286730 75134
rect 286966 74898 287008 75134
rect 286688 74866 287008 74898
rect 317408 75454 317728 75486
rect 317408 75218 317450 75454
rect 317686 75218 317728 75454
rect 317408 75134 317728 75218
rect 317408 74898 317450 75134
rect 317686 74898 317728 75134
rect 317408 74866 317728 74898
rect 348128 75454 348448 75486
rect 348128 75218 348170 75454
rect 348406 75218 348448 75454
rect 348128 75134 348448 75218
rect 348128 74898 348170 75134
rect 348406 74898 348448 75134
rect 348128 74866 348448 74898
rect 378848 75454 379168 75486
rect 378848 75218 378890 75454
rect 379126 75218 379168 75454
rect 378848 75134 379168 75218
rect 378848 74898 378890 75134
rect 379126 74898 379168 75134
rect 378848 74866 379168 74898
rect 409568 75454 409888 75486
rect 409568 75218 409610 75454
rect 409846 75218 409888 75454
rect 409568 75134 409888 75218
rect 409568 74898 409610 75134
rect 409846 74898 409888 75134
rect 409568 74866 409888 74898
rect 440288 75454 440608 75486
rect 440288 75218 440330 75454
rect 440566 75218 440608 75454
rect 440288 75134 440608 75218
rect 440288 74898 440330 75134
rect 440566 74898 440608 75134
rect 440288 74866 440608 74898
rect 471008 75454 471328 75486
rect 471008 75218 471050 75454
rect 471286 75218 471328 75454
rect 471008 75134 471328 75218
rect 471008 74898 471050 75134
rect 471286 74898 471328 75134
rect 471008 74866 471328 74898
rect 501728 75454 502048 75486
rect 501728 75218 501770 75454
rect 502006 75218 502048 75454
rect 501728 75134 502048 75218
rect 501728 74898 501770 75134
rect 502006 74898 502048 75134
rect 501728 74866 502048 74898
rect 532448 75454 532768 75486
rect 532448 75218 532490 75454
rect 532726 75218 532768 75454
rect 532448 75134 532768 75218
rect 532448 74898 532490 75134
rect 532726 74898 532768 75134
rect 532448 74866 532768 74898
rect 563168 75454 563488 75486
rect 563168 75218 563210 75454
rect 563446 75218 563488 75454
rect 563168 75134 563488 75218
rect 563168 74898 563210 75134
rect 563446 74898 563488 75134
rect 563168 74866 563488 74898
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 25568 43174 25888 43206
rect 25568 42938 25610 43174
rect 25846 42938 25888 43174
rect 25568 42854 25888 42938
rect 25568 42618 25610 42854
rect 25846 42618 25888 42854
rect 25568 42586 25888 42618
rect 56288 43174 56608 43206
rect 56288 42938 56330 43174
rect 56566 42938 56608 43174
rect 56288 42854 56608 42938
rect 56288 42618 56330 42854
rect 56566 42618 56608 42854
rect 56288 42586 56608 42618
rect 87008 43174 87328 43206
rect 87008 42938 87050 43174
rect 87286 42938 87328 43174
rect 87008 42854 87328 42938
rect 87008 42618 87050 42854
rect 87286 42618 87328 42854
rect 87008 42586 87328 42618
rect 117728 43174 118048 43206
rect 117728 42938 117770 43174
rect 118006 42938 118048 43174
rect 117728 42854 118048 42938
rect 117728 42618 117770 42854
rect 118006 42618 118048 42854
rect 117728 42586 118048 42618
rect 148448 43174 148768 43206
rect 148448 42938 148490 43174
rect 148726 42938 148768 43174
rect 148448 42854 148768 42938
rect 148448 42618 148490 42854
rect 148726 42618 148768 42854
rect 148448 42586 148768 42618
rect 179168 43174 179488 43206
rect 179168 42938 179210 43174
rect 179446 42938 179488 43174
rect 179168 42854 179488 42938
rect 179168 42618 179210 42854
rect 179446 42618 179488 42854
rect 179168 42586 179488 42618
rect 209888 43174 210208 43206
rect 209888 42938 209930 43174
rect 210166 42938 210208 43174
rect 209888 42854 210208 42938
rect 209888 42618 209930 42854
rect 210166 42618 210208 42854
rect 209888 42586 210208 42618
rect 240608 43174 240928 43206
rect 240608 42938 240650 43174
rect 240886 42938 240928 43174
rect 240608 42854 240928 42938
rect 240608 42618 240650 42854
rect 240886 42618 240928 42854
rect 240608 42586 240928 42618
rect 271328 43174 271648 43206
rect 271328 42938 271370 43174
rect 271606 42938 271648 43174
rect 271328 42854 271648 42938
rect 271328 42618 271370 42854
rect 271606 42618 271648 42854
rect 271328 42586 271648 42618
rect 302048 43174 302368 43206
rect 302048 42938 302090 43174
rect 302326 42938 302368 43174
rect 302048 42854 302368 42938
rect 302048 42618 302090 42854
rect 302326 42618 302368 42854
rect 302048 42586 302368 42618
rect 332768 43174 333088 43206
rect 332768 42938 332810 43174
rect 333046 42938 333088 43174
rect 332768 42854 333088 42938
rect 332768 42618 332810 42854
rect 333046 42618 333088 42854
rect 332768 42586 333088 42618
rect 363488 43174 363808 43206
rect 363488 42938 363530 43174
rect 363766 42938 363808 43174
rect 363488 42854 363808 42938
rect 363488 42618 363530 42854
rect 363766 42618 363808 42854
rect 363488 42586 363808 42618
rect 394208 43174 394528 43206
rect 394208 42938 394250 43174
rect 394486 42938 394528 43174
rect 394208 42854 394528 42938
rect 394208 42618 394250 42854
rect 394486 42618 394528 42854
rect 394208 42586 394528 42618
rect 424928 43174 425248 43206
rect 424928 42938 424970 43174
rect 425206 42938 425248 43174
rect 424928 42854 425248 42938
rect 424928 42618 424970 42854
rect 425206 42618 425248 42854
rect 424928 42586 425248 42618
rect 455648 43174 455968 43206
rect 455648 42938 455690 43174
rect 455926 42938 455968 43174
rect 455648 42854 455968 42938
rect 455648 42618 455690 42854
rect 455926 42618 455968 42854
rect 455648 42586 455968 42618
rect 486368 43174 486688 43206
rect 486368 42938 486410 43174
rect 486646 42938 486688 43174
rect 486368 42854 486688 42938
rect 486368 42618 486410 42854
rect 486646 42618 486688 42854
rect 486368 42586 486688 42618
rect 517088 43174 517408 43206
rect 517088 42938 517130 43174
rect 517366 42938 517408 43174
rect 517088 42854 517408 42938
rect 517088 42618 517130 42854
rect 517366 42618 517408 42854
rect 517088 42586 517408 42618
rect 547808 43174 548128 43206
rect 547808 42938 547850 43174
rect 548086 42938 548128 43174
rect 547808 42854 548128 42938
rect 547808 42618 547850 42854
rect 548086 42618 548128 42854
rect 547808 42586 548128 42618
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 10208 39454 10528 39486
rect 10208 39218 10250 39454
rect 10486 39218 10528 39454
rect 10208 39134 10528 39218
rect 10208 38898 10250 39134
rect 10486 38898 10528 39134
rect 10208 38866 10528 38898
rect 40928 39454 41248 39486
rect 40928 39218 40970 39454
rect 41206 39218 41248 39454
rect 40928 39134 41248 39218
rect 40928 38898 40970 39134
rect 41206 38898 41248 39134
rect 40928 38866 41248 38898
rect 71648 39454 71968 39486
rect 71648 39218 71690 39454
rect 71926 39218 71968 39454
rect 71648 39134 71968 39218
rect 71648 38898 71690 39134
rect 71926 38898 71968 39134
rect 71648 38866 71968 38898
rect 102368 39454 102688 39486
rect 102368 39218 102410 39454
rect 102646 39218 102688 39454
rect 102368 39134 102688 39218
rect 102368 38898 102410 39134
rect 102646 38898 102688 39134
rect 102368 38866 102688 38898
rect 133088 39454 133408 39486
rect 133088 39218 133130 39454
rect 133366 39218 133408 39454
rect 133088 39134 133408 39218
rect 133088 38898 133130 39134
rect 133366 38898 133408 39134
rect 133088 38866 133408 38898
rect 163808 39454 164128 39486
rect 163808 39218 163850 39454
rect 164086 39218 164128 39454
rect 163808 39134 164128 39218
rect 163808 38898 163850 39134
rect 164086 38898 164128 39134
rect 163808 38866 164128 38898
rect 194528 39454 194848 39486
rect 194528 39218 194570 39454
rect 194806 39218 194848 39454
rect 194528 39134 194848 39218
rect 194528 38898 194570 39134
rect 194806 38898 194848 39134
rect 194528 38866 194848 38898
rect 225248 39454 225568 39486
rect 225248 39218 225290 39454
rect 225526 39218 225568 39454
rect 225248 39134 225568 39218
rect 225248 38898 225290 39134
rect 225526 38898 225568 39134
rect 225248 38866 225568 38898
rect 255968 39454 256288 39486
rect 255968 39218 256010 39454
rect 256246 39218 256288 39454
rect 255968 39134 256288 39218
rect 255968 38898 256010 39134
rect 256246 38898 256288 39134
rect 255968 38866 256288 38898
rect 286688 39454 287008 39486
rect 286688 39218 286730 39454
rect 286966 39218 287008 39454
rect 286688 39134 287008 39218
rect 286688 38898 286730 39134
rect 286966 38898 287008 39134
rect 286688 38866 287008 38898
rect 317408 39454 317728 39486
rect 317408 39218 317450 39454
rect 317686 39218 317728 39454
rect 317408 39134 317728 39218
rect 317408 38898 317450 39134
rect 317686 38898 317728 39134
rect 317408 38866 317728 38898
rect 348128 39454 348448 39486
rect 348128 39218 348170 39454
rect 348406 39218 348448 39454
rect 348128 39134 348448 39218
rect 348128 38898 348170 39134
rect 348406 38898 348448 39134
rect 348128 38866 348448 38898
rect 378848 39454 379168 39486
rect 378848 39218 378890 39454
rect 379126 39218 379168 39454
rect 378848 39134 379168 39218
rect 378848 38898 378890 39134
rect 379126 38898 379168 39134
rect 378848 38866 379168 38898
rect 409568 39454 409888 39486
rect 409568 39218 409610 39454
rect 409846 39218 409888 39454
rect 409568 39134 409888 39218
rect 409568 38898 409610 39134
rect 409846 38898 409888 39134
rect 409568 38866 409888 38898
rect 440288 39454 440608 39486
rect 440288 39218 440330 39454
rect 440566 39218 440608 39454
rect 440288 39134 440608 39218
rect 440288 38898 440330 39134
rect 440566 38898 440608 39134
rect 440288 38866 440608 38898
rect 471008 39454 471328 39486
rect 471008 39218 471050 39454
rect 471286 39218 471328 39454
rect 471008 39134 471328 39218
rect 471008 38898 471050 39134
rect 471286 38898 471328 39134
rect 471008 38866 471328 38898
rect 501728 39454 502048 39486
rect 501728 39218 501770 39454
rect 502006 39218 502048 39454
rect 501728 39134 502048 39218
rect 501728 38898 501770 39134
rect 502006 38898 502048 39134
rect 501728 38866 502048 38898
rect 532448 39454 532768 39486
rect 532448 39218 532490 39454
rect 532726 39218 532768 39454
rect 532448 39134 532768 39218
rect 532448 38898 532490 39134
rect 532726 38898 532768 39134
rect 532448 38866 532768 38898
rect 563168 39454 563488 39486
rect 563168 39218 563210 39454
rect 563446 39218 563488 39454
rect 563168 39134 563488 39218
rect 563168 38898 563210 39134
rect 563446 38898 563488 39134
rect 563168 38866 563488 38898
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 5514 7174 6134 7375
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect 5514 -1306 6134 6618
rect 5514 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 6134 -1306
rect 5514 -1626 6134 -1542
rect 5514 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 6134 -1626
rect 5514 -7654 6134 -1862
rect 37794 3454 38414 7375
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 41514 7174 42134 7375
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -1306 42134 6618
rect 41514 -1542 41546 -1306
rect 41782 -1542 41866 -1306
rect 42102 -1542 42134 -1306
rect 41514 -1626 42134 -1542
rect 41514 -1862 41546 -1626
rect 41782 -1862 41866 -1626
rect 42102 -1862 42134 -1626
rect 41514 -7654 42134 -1862
rect 73794 3454 74414 7375
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 77514 7174 78134 7375
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -1306 78134 6618
rect 77514 -1542 77546 -1306
rect 77782 -1542 77866 -1306
rect 78102 -1542 78134 -1306
rect 77514 -1626 78134 -1542
rect 77514 -1862 77546 -1626
rect 77782 -1862 77866 -1626
rect 78102 -1862 78134 -1626
rect 77514 -7654 78134 -1862
rect 109794 3454 110414 7375
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 113514 7174 114134 7375
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -1306 114134 6618
rect 113514 -1542 113546 -1306
rect 113782 -1542 113866 -1306
rect 114102 -1542 114134 -1306
rect 113514 -1626 114134 -1542
rect 113514 -1862 113546 -1626
rect 113782 -1862 113866 -1626
rect 114102 -1862 114134 -1626
rect 113514 -7654 114134 -1862
rect 145794 3454 146414 7375
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 149514 7174 150134 7375
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -1306 150134 6618
rect 149514 -1542 149546 -1306
rect 149782 -1542 149866 -1306
rect 150102 -1542 150134 -1306
rect 149514 -1626 150134 -1542
rect 149514 -1862 149546 -1626
rect 149782 -1862 149866 -1626
rect 150102 -1862 150134 -1626
rect 149514 -7654 150134 -1862
rect 181794 3454 182414 7375
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 185514 7174 186134 7375
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -1306 186134 6618
rect 185514 -1542 185546 -1306
rect 185782 -1542 185866 -1306
rect 186102 -1542 186134 -1306
rect 185514 -1626 186134 -1542
rect 185514 -1862 185546 -1626
rect 185782 -1862 185866 -1626
rect 186102 -1862 186134 -1626
rect 185514 -7654 186134 -1862
rect 217794 3454 218414 7375
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 221514 7174 222134 7375
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -1306 222134 6618
rect 221514 -1542 221546 -1306
rect 221782 -1542 221866 -1306
rect 222102 -1542 222134 -1306
rect 221514 -1626 222134 -1542
rect 221514 -1862 221546 -1626
rect 221782 -1862 221866 -1626
rect 222102 -1862 222134 -1626
rect 221514 -7654 222134 -1862
rect 253794 3454 254414 7375
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 257514 7174 258134 7375
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -1306 258134 6618
rect 257514 -1542 257546 -1306
rect 257782 -1542 257866 -1306
rect 258102 -1542 258134 -1306
rect 257514 -1626 258134 -1542
rect 257514 -1862 257546 -1626
rect 257782 -1862 257866 -1626
rect 258102 -1862 258134 -1626
rect 257514 -7654 258134 -1862
rect 289794 3454 290414 7375
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 293514 7174 294134 7375
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -1306 294134 6618
rect 293514 -1542 293546 -1306
rect 293782 -1542 293866 -1306
rect 294102 -1542 294134 -1306
rect 293514 -1626 294134 -1542
rect 293514 -1862 293546 -1626
rect 293782 -1862 293866 -1626
rect 294102 -1862 294134 -1626
rect 293514 -7654 294134 -1862
rect 325794 3454 326414 7375
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 329514 7174 330134 7375
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -1306 330134 6618
rect 329514 -1542 329546 -1306
rect 329782 -1542 329866 -1306
rect 330102 -1542 330134 -1306
rect 329514 -1626 330134 -1542
rect 329514 -1862 329546 -1626
rect 329782 -1862 329866 -1626
rect 330102 -1862 330134 -1626
rect 329514 -7654 330134 -1862
rect 361794 3454 362414 7375
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 365514 7174 366134 7375
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -1306 366134 6618
rect 365514 -1542 365546 -1306
rect 365782 -1542 365866 -1306
rect 366102 -1542 366134 -1306
rect 365514 -1626 366134 -1542
rect 365514 -1862 365546 -1626
rect 365782 -1862 365866 -1626
rect 366102 -1862 366134 -1626
rect 365514 -7654 366134 -1862
rect 397794 3454 398414 7375
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 401514 7174 402134 7375
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -1306 402134 6618
rect 401514 -1542 401546 -1306
rect 401782 -1542 401866 -1306
rect 402102 -1542 402134 -1306
rect 401514 -1626 402134 -1542
rect 401514 -1862 401546 -1626
rect 401782 -1862 401866 -1626
rect 402102 -1862 402134 -1626
rect 401514 -7654 402134 -1862
rect 433794 3454 434414 7375
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 437514 7174 438134 7375
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -1306 438134 6618
rect 437514 -1542 437546 -1306
rect 437782 -1542 437866 -1306
rect 438102 -1542 438134 -1306
rect 437514 -1626 438134 -1542
rect 437514 -1862 437546 -1626
rect 437782 -1862 437866 -1626
rect 438102 -1862 438134 -1626
rect 437514 -7654 438134 -1862
rect 469794 3454 470414 7375
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 473514 7174 474134 7375
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -1306 474134 6618
rect 473514 -1542 473546 -1306
rect 473782 -1542 473866 -1306
rect 474102 -1542 474134 -1306
rect 473514 -1626 474134 -1542
rect 473514 -1862 473546 -1626
rect 473782 -1862 473866 -1626
rect 474102 -1862 474134 -1626
rect 473514 -7654 474134 -1862
rect 505794 3454 506414 7375
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 509514 7174 510134 7375
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -1306 510134 6618
rect 509514 -1542 509546 -1306
rect 509782 -1542 509866 -1306
rect 510102 -1542 510134 -1306
rect 509514 -1626 510134 -1542
rect 509514 -1862 509546 -1626
rect 509782 -1862 509866 -1626
rect 510102 -1862 510134 -1626
rect 509514 -7654 510134 -1862
rect 541794 3454 542414 7375
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 545514 7174 546134 7375
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -1306 546134 6618
rect 545514 -1542 545546 -1306
rect 545782 -1542 545866 -1306
rect 546102 -1542 546134 -1306
rect 545514 -1626 546134 -1542
rect 545514 -1862 545546 -1626
rect 545782 -1862 545866 -1626
rect 546102 -1862 546134 -1626
rect 545514 -7654 546134 -1862
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 581514 705798 582134 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 581514 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 582134 705798
rect 581514 705478 582134 705562
rect 581514 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 582134 705478
rect 581514 691174 582134 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -1306 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691174 586890 705242
rect 586270 690938 586302 691174
rect 586538 690938 586622 691174
rect 586858 690938 586890 691174
rect 586270 690854 586890 690938
rect 586270 690618 586302 690854
rect 586538 690618 586622 690854
rect 586858 690618 586890 690854
rect 586270 655174 586890 690618
rect 586270 654938 586302 655174
rect 586538 654938 586622 655174
rect 586858 654938 586890 655174
rect 586270 654854 586890 654938
rect 586270 654618 586302 654854
rect 586538 654618 586622 654854
rect 586858 654618 586890 654854
rect 586270 619174 586890 654618
rect 586270 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 586890 619174
rect 586270 618854 586890 618938
rect 586270 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 586890 618854
rect 586270 583174 586890 618618
rect 586270 582938 586302 583174
rect 586538 582938 586622 583174
rect 586858 582938 586890 583174
rect 586270 582854 586890 582938
rect 586270 582618 586302 582854
rect 586538 582618 586622 582854
rect 586858 582618 586890 582854
rect 586270 547174 586890 582618
rect 586270 546938 586302 547174
rect 586538 546938 586622 547174
rect 586858 546938 586890 547174
rect 586270 546854 586890 546938
rect 586270 546618 586302 546854
rect 586538 546618 586622 546854
rect 586858 546618 586890 546854
rect 586270 511174 586890 546618
rect 586270 510938 586302 511174
rect 586538 510938 586622 511174
rect 586858 510938 586890 511174
rect 586270 510854 586890 510938
rect 586270 510618 586302 510854
rect 586538 510618 586622 510854
rect 586858 510618 586890 510854
rect 586270 475174 586890 510618
rect 586270 474938 586302 475174
rect 586538 474938 586622 475174
rect 586858 474938 586890 475174
rect 586270 474854 586890 474938
rect 586270 474618 586302 474854
rect 586538 474618 586622 474854
rect 586858 474618 586890 474854
rect 586270 439174 586890 474618
rect 586270 438938 586302 439174
rect 586538 438938 586622 439174
rect 586858 438938 586890 439174
rect 586270 438854 586890 438938
rect 586270 438618 586302 438854
rect 586538 438618 586622 438854
rect 586858 438618 586890 438854
rect 586270 403174 586890 438618
rect 586270 402938 586302 403174
rect 586538 402938 586622 403174
rect 586858 402938 586890 403174
rect 586270 402854 586890 402938
rect 586270 402618 586302 402854
rect 586538 402618 586622 402854
rect 586858 402618 586890 402854
rect 586270 367174 586890 402618
rect 586270 366938 586302 367174
rect 586538 366938 586622 367174
rect 586858 366938 586890 367174
rect 586270 366854 586890 366938
rect 586270 366618 586302 366854
rect 586538 366618 586622 366854
rect 586858 366618 586890 366854
rect 586270 331174 586890 366618
rect 586270 330938 586302 331174
rect 586538 330938 586622 331174
rect 586858 330938 586890 331174
rect 586270 330854 586890 330938
rect 586270 330618 586302 330854
rect 586538 330618 586622 330854
rect 586858 330618 586890 330854
rect 586270 295174 586890 330618
rect 586270 294938 586302 295174
rect 586538 294938 586622 295174
rect 586858 294938 586890 295174
rect 586270 294854 586890 294938
rect 586270 294618 586302 294854
rect 586538 294618 586622 294854
rect 586858 294618 586890 294854
rect 586270 259174 586890 294618
rect 586270 258938 586302 259174
rect 586538 258938 586622 259174
rect 586858 258938 586890 259174
rect 586270 258854 586890 258938
rect 586270 258618 586302 258854
rect 586538 258618 586622 258854
rect 586858 258618 586890 258854
rect 586270 223174 586890 258618
rect 586270 222938 586302 223174
rect 586538 222938 586622 223174
rect 586858 222938 586890 223174
rect 586270 222854 586890 222938
rect 586270 222618 586302 222854
rect 586538 222618 586622 222854
rect 586858 222618 586890 222854
rect 586270 187174 586890 222618
rect 586270 186938 586302 187174
rect 586538 186938 586622 187174
rect 586858 186938 586890 187174
rect 586270 186854 586890 186938
rect 586270 186618 586302 186854
rect 586538 186618 586622 186854
rect 586858 186618 586890 186854
rect 586270 151174 586890 186618
rect 586270 150938 586302 151174
rect 586538 150938 586622 151174
rect 586858 150938 586890 151174
rect 586270 150854 586890 150938
rect 586270 150618 586302 150854
rect 586538 150618 586622 150854
rect 586858 150618 586890 150854
rect 586270 115174 586890 150618
rect 586270 114938 586302 115174
rect 586538 114938 586622 115174
rect 586858 114938 586890 115174
rect 586270 114854 586890 114938
rect 586270 114618 586302 114854
rect 586538 114618 586622 114854
rect 586858 114618 586890 114854
rect 586270 79174 586890 114618
rect 586270 78938 586302 79174
rect 586538 78938 586622 79174
rect 586858 78938 586890 79174
rect 586270 78854 586890 78938
rect 586270 78618 586302 78854
rect 586538 78618 586622 78854
rect 586858 78618 586890 78854
rect 586270 43174 586890 78618
rect 586270 42938 586302 43174
rect 586538 42938 586622 43174
rect 586858 42938 586890 43174
rect 586270 42854 586890 42938
rect 586270 42618 586302 42854
rect 586538 42618 586622 42854
rect 586858 42618 586890 42854
rect 586270 7174 586890 42618
rect 586270 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 586890 7174
rect 586270 6854 586890 6938
rect 586270 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 586890 6854
rect 581514 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 582134 -1306
rect 581514 -1626 582134 -1542
rect 581514 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 582134 -1626
rect 581514 -7654 582134 -1862
rect 586270 -1306 586890 6618
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 694894 587850 706202
rect 587230 694658 587262 694894
rect 587498 694658 587582 694894
rect 587818 694658 587850 694894
rect 587230 694574 587850 694658
rect 587230 694338 587262 694574
rect 587498 694338 587582 694574
rect 587818 694338 587850 694574
rect 587230 658894 587850 694338
rect 587230 658658 587262 658894
rect 587498 658658 587582 658894
rect 587818 658658 587850 658894
rect 587230 658574 587850 658658
rect 587230 658338 587262 658574
rect 587498 658338 587582 658574
rect 587818 658338 587850 658574
rect 587230 622894 587850 658338
rect 587230 622658 587262 622894
rect 587498 622658 587582 622894
rect 587818 622658 587850 622894
rect 587230 622574 587850 622658
rect 587230 622338 587262 622574
rect 587498 622338 587582 622574
rect 587818 622338 587850 622574
rect 587230 586894 587850 622338
rect 587230 586658 587262 586894
rect 587498 586658 587582 586894
rect 587818 586658 587850 586894
rect 587230 586574 587850 586658
rect 587230 586338 587262 586574
rect 587498 586338 587582 586574
rect 587818 586338 587850 586574
rect 587230 550894 587850 586338
rect 587230 550658 587262 550894
rect 587498 550658 587582 550894
rect 587818 550658 587850 550894
rect 587230 550574 587850 550658
rect 587230 550338 587262 550574
rect 587498 550338 587582 550574
rect 587818 550338 587850 550574
rect 587230 514894 587850 550338
rect 587230 514658 587262 514894
rect 587498 514658 587582 514894
rect 587818 514658 587850 514894
rect 587230 514574 587850 514658
rect 587230 514338 587262 514574
rect 587498 514338 587582 514574
rect 587818 514338 587850 514574
rect 587230 478894 587850 514338
rect 587230 478658 587262 478894
rect 587498 478658 587582 478894
rect 587818 478658 587850 478894
rect 587230 478574 587850 478658
rect 587230 478338 587262 478574
rect 587498 478338 587582 478574
rect 587818 478338 587850 478574
rect 587230 442894 587850 478338
rect 587230 442658 587262 442894
rect 587498 442658 587582 442894
rect 587818 442658 587850 442894
rect 587230 442574 587850 442658
rect 587230 442338 587262 442574
rect 587498 442338 587582 442574
rect 587818 442338 587850 442574
rect 587230 406894 587850 442338
rect 587230 406658 587262 406894
rect 587498 406658 587582 406894
rect 587818 406658 587850 406894
rect 587230 406574 587850 406658
rect 587230 406338 587262 406574
rect 587498 406338 587582 406574
rect 587818 406338 587850 406574
rect 587230 370894 587850 406338
rect 587230 370658 587262 370894
rect 587498 370658 587582 370894
rect 587818 370658 587850 370894
rect 587230 370574 587850 370658
rect 587230 370338 587262 370574
rect 587498 370338 587582 370574
rect 587818 370338 587850 370574
rect 587230 334894 587850 370338
rect 587230 334658 587262 334894
rect 587498 334658 587582 334894
rect 587818 334658 587850 334894
rect 587230 334574 587850 334658
rect 587230 334338 587262 334574
rect 587498 334338 587582 334574
rect 587818 334338 587850 334574
rect 587230 298894 587850 334338
rect 587230 298658 587262 298894
rect 587498 298658 587582 298894
rect 587818 298658 587850 298894
rect 587230 298574 587850 298658
rect 587230 298338 587262 298574
rect 587498 298338 587582 298574
rect 587818 298338 587850 298574
rect 587230 262894 587850 298338
rect 587230 262658 587262 262894
rect 587498 262658 587582 262894
rect 587818 262658 587850 262894
rect 587230 262574 587850 262658
rect 587230 262338 587262 262574
rect 587498 262338 587582 262574
rect 587818 262338 587850 262574
rect 587230 226894 587850 262338
rect 587230 226658 587262 226894
rect 587498 226658 587582 226894
rect 587818 226658 587850 226894
rect 587230 226574 587850 226658
rect 587230 226338 587262 226574
rect 587498 226338 587582 226574
rect 587818 226338 587850 226574
rect 587230 190894 587850 226338
rect 587230 190658 587262 190894
rect 587498 190658 587582 190894
rect 587818 190658 587850 190894
rect 587230 190574 587850 190658
rect 587230 190338 587262 190574
rect 587498 190338 587582 190574
rect 587818 190338 587850 190574
rect 587230 154894 587850 190338
rect 587230 154658 587262 154894
rect 587498 154658 587582 154894
rect 587818 154658 587850 154894
rect 587230 154574 587850 154658
rect 587230 154338 587262 154574
rect 587498 154338 587582 154574
rect 587818 154338 587850 154574
rect 587230 118894 587850 154338
rect 587230 118658 587262 118894
rect 587498 118658 587582 118894
rect 587818 118658 587850 118894
rect 587230 118574 587850 118658
rect 587230 118338 587262 118574
rect 587498 118338 587582 118574
rect 587818 118338 587850 118574
rect 587230 82894 587850 118338
rect 587230 82658 587262 82894
rect 587498 82658 587582 82894
rect 587818 82658 587850 82894
rect 587230 82574 587850 82658
rect 587230 82338 587262 82574
rect 587498 82338 587582 82574
rect 587818 82338 587850 82574
rect 587230 46894 587850 82338
rect 587230 46658 587262 46894
rect 587498 46658 587582 46894
rect 587818 46658 587850 46894
rect 587230 46574 587850 46658
rect 587230 46338 587262 46574
rect 587498 46338 587582 46574
rect 587818 46338 587850 46574
rect 587230 10894 587850 46338
rect 587230 10658 587262 10894
rect 587498 10658 587582 10894
rect 587818 10658 587850 10894
rect 587230 10574 587850 10658
rect 587230 10338 587262 10574
rect 587498 10338 587582 10574
rect 587818 10338 587850 10574
rect 587230 -2266 587850 10338
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 698614 588810 707162
rect 588190 698378 588222 698614
rect 588458 698378 588542 698614
rect 588778 698378 588810 698614
rect 588190 698294 588810 698378
rect 588190 698058 588222 698294
rect 588458 698058 588542 698294
rect 588778 698058 588810 698294
rect 588190 662614 588810 698058
rect 588190 662378 588222 662614
rect 588458 662378 588542 662614
rect 588778 662378 588810 662614
rect 588190 662294 588810 662378
rect 588190 662058 588222 662294
rect 588458 662058 588542 662294
rect 588778 662058 588810 662294
rect 588190 626614 588810 662058
rect 588190 626378 588222 626614
rect 588458 626378 588542 626614
rect 588778 626378 588810 626614
rect 588190 626294 588810 626378
rect 588190 626058 588222 626294
rect 588458 626058 588542 626294
rect 588778 626058 588810 626294
rect 588190 590614 588810 626058
rect 588190 590378 588222 590614
rect 588458 590378 588542 590614
rect 588778 590378 588810 590614
rect 588190 590294 588810 590378
rect 588190 590058 588222 590294
rect 588458 590058 588542 590294
rect 588778 590058 588810 590294
rect 588190 554614 588810 590058
rect 588190 554378 588222 554614
rect 588458 554378 588542 554614
rect 588778 554378 588810 554614
rect 588190 554294 588810 554378
rect 588190 554058 588222 554294
rect 588458 554058 588542 554294
rect 588778 554058 588810 554294
rect 588190 518614 588810 554058
rect 588190 518378 588222 518614
rect 588458 518378 588542 518614
rect 588778 518378 588810 518614
rect 588190 518294 588810 518378
rect 588190 518058 588222 518294
rect 588458 518058 588542 518294
rect 588778 518058 588810 518294
rect 588190 482614 588810 518058
rect 588190 482378 588222 482614
rect 588458 482378 588542 482614
rect 588778 482378 588810 482614
rect 588190 482294 588810 482378
rect 588190 482058 588222 482294
rect 588458 482058 588542 482294
rect 588778 482058 588810 482294
rect 588190 446614 588810 482058
rect 588190 446378 588222 446614
rect 588458 446378 588542 446614
rect 588778 446378 588810 446614
rect 588190 446294 588810 446378
rect 588190 446058 588222 446294
rect 588458 446058 588542 446294
rect 588778 446058 588810 446294
rect 588190 410614 588810 446058
rect 588190 410378 588222 410614
rect 588458 410378 588542 410614
rect 588778 410378 588810 410614
rect 588190 410294 588810 410378
rect 588190 410058 588222 410294
rect 588458 410058 588542 410294
rect 588778 410058 588810 410294
rect 588190 374614 588810 410058
rect 588190 374378 588222 374614
rect 588458 374378 588542 374614
rect 588778 374378 588810 374614
rect 588190 374294 588810 374378
rect 588190 374058 588222 374294
rect 588458 374058 588542 374294
rect 588778 374058 588810 374294
rect 588190 338614 588810 374058
rect 588190 338378 588222 338614
rect 588458 338378 588542 338614
rect 588778 338378 588810 338614
rect 588190 338294 588810 338378
rect 588190 338058 588222 338294
rect 588458 338058 588542 338294
rect 588778 338058 588810 338294
rect 588190 302614 588810 338058
rect 588190 302378 588222 302614
rect 588458 302378 588542 302614
rect 588778 302378 588810 302614
rect 588190 302294 588810 302378
rect 588190 302058 588222 302294
rect 588458 302058 588542 302294
rect 588778 302058 588810 302294
rect 588190 266614 588810 302058
rect 588190 266378 588222 266614
rect 588458 266378 588542 266614
rect 588778 266378 588810 266614
rect 588190 266294 588810 266378
rect 588190 266058 588222 266294
rect 588458 266058 588542 266294
rect 588778 266058 588810 266294
rect 588190 230614 588810 266058
rect 588190 230378 588222 230614
rect 588458 230378 588542 230614
rect 588778 230378 588810 230614
rect 588190 230294 588810 230378
rect 588190 230058 588222 230294
rect 588458 230058 588542 230294
rect 588778 230058 588810 230294
rect 588190 194614 588810 230058
rect 588190 194378 588222 194614
rect 588458 194378 588542 194614
rect 588778 194378 588810 194614
rect 588190 194294 588810 194378
rect 588190 194058 588222 194294
rect 588458 194058 588542 194294
rect 588778 194058 588810 194294
rect 588190 158614 588810 194058
rect 588190 158378 588222 158614
rect 588458 158378 588542 158614
rect 588778 158378 588810 158614
rect 588190 158294 588810 158378
rect 588190 158058 588222 158294
rect 588458 158058 588542 158294
rect 588778 158058 588810 158294
rect 588190 122614 588810 158058
rect 588190 122378 588222 122614
rect 588458 122378 588542 122614
rect 588778 122378 588810 122614
rect 588190 122294 588810 122378
rect 588190 122058 588222 122294
rect 588458 122058 588542 122294
rect 588778 122058 588810 122294
rect 588190 86614 588810 122058
rect 588190 86378 588222 86614
rect 588458 86378 588542 86614
rect 588778 86378 588810 86614
rect 588190 86294 588810 86378
rect 588190 86058 588222 86294
rect 588458 86058 588542 86294
rect 588778 86058 588810 86294
rect 588190 50614 588810 86058
rect 588190 50378 588222 50614
rect 588458 50378 588542 50614
rect 588778 50378 588810 50614
rect 588190 50294 588810 50378
rect 588190 50058 588222 50294
rect 588458 50058 588542 50294
rect 588778 50058 588810 50294
rect 588190 14614 588810 50058
rect 588190 14378 588222 14614
rect 588458 14378 588542 14614
rect 588778 14378 588810 14614
rect 588190 14294 588810 14378
rect 588190 14058 588222 14294
rect 588458 14058 588542 14294
rect 588778 14058 588810 14294
rect 588190 -3226 588810 14058
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 666334 589770 708122
rect 589150 666098 589182 666334
rect 589418 666098 589502 666334
rect 589738 666098 589770 666334
rect 589150 666014 589770 666098
rect 589150 665778 589182 666014
rect 589418 665778 589502 666014
rect 589738 665778 589770 666014
rect 589150 630334 589770 665778
rect 589150 630098 589182 630334
rect 589418 630098 589502 630334
rect 589738 630098 589770 630334
rect 589150 630014 589770 630098
rect 589150 629778 589182 630014
rect 589418 629778 589502 630014
rect 589738 629778 589770 630014
rect 589150 594334 589770 629778
rect 589150 594098 589182 594334
rect 589418 594098 589502 594334
rect 589738 594098 589770 594334
rect 589150 594014 589770 594098
rect 589150 593778 589182 594014
rect 589418 593778 589502 594014
rect 589738 593778 589770 594014
rect 589150 558334 589770 593778
rect 589150 558098 589182 558334
rect 589418 558098 589502 558334
rect 589738 558098 589770 558334
rect 589150 558014 589770 558098
rect 589150 557778 589182 558014
rect 589418 557778 589502 558014
rect 589738 557778 589770 558014
rect 589150 522334 589770 557778
rect 589150 522098 589182 522334
rect 589418 522098 589502 522334
rect 589738 522098 589770 522334
rect 589150 522014 589770 522098
rect 589150 521778 589182 522014
rect 589418 521778 589502 522014
rect 589738 521778 589770 522014
rect 589150 486334 589770 521778
rect 589150 486098 589182 486334
rect 589418 486098 589502 486334
rect 589738 486098 589770 486334
rect 589150 486014 589770 486098
rect 589150 485778 589182 486014
rect 589418 485778 589502 486014
rect 589738 485778 589770 486014
rect 589150 450334 589770 485778
rect 589150 450098 589182 450334
rect 589418 450098 589502 450334
rect 589738 450098 589770 450334
rect 589150 450014 589770 450098
rect 589150 449778 589182 450014
rect 589418 449778 589502 450014
rect 589738 449778 589770 450014
rect 589150 414334 589770 449778
rect 589150 414098 589182 414334
rect 589418 414098 589502 414334
rect 589738 414098 589770 414334
rect 589150 414014 589770 414098
rect 589150 413778 589182 414014
rect 589418 413778 589502 414014
rect 589738 413778 589770 414014
rect 589150 378334 589770 413778
rect 589150 378098 589182 378334
rect 589418 378098 589502 378334
rect 589738 378098 589770 378334
rect 589150 378014 589770 378098
rect 589150 377778 589182 378014
rect 589418 377778 589502 378014
rect 589738 377778 589770 378014
rect 589150 342334 589770 377778
rect 589150 342098 589182 342334
rect 589418 342098 589502 342334
rect 589738 342098 589770 342334
rect 589150 342014 589770 342098
rect 589150 341778 589182 342014
rect 589418 341778 589502 342014
rect 589738 341778 589770 342014
rect 589150 306334 589770 341778
rect 589150 306098 589182 306334
rect 589418 306098 589502 306334
rect 589738 306098 589770 306334
rect 589150 306014 589770 306098
rect 589150 305778 589182 306014
rect 589418 305778 589502 306014
rect 589738 305778 589770 306014
rect 589150 270334 589770 305778
rect 589150 270098 589182 270334
rect 589418 270098 589502 270334
rect 589738 270098 589770 270334
rect 589150 270014 589770 270098
rect 589150 269778 589182 270014
rect 589418 269778 589502 270014
rect 589738 269778 589770 270014
rect 589150 234334 589770 269778
rect 589150 234098 589182 234334
rect 589418 234098 589502 234334
rect 589738 234098 589770 234334
rect 589150 234014 589770 234098
rect 589150 233778 589182 234014
rect 589418 233778 589502 234014
rect 589738 233778 589770 234014
rect 589150 198334 589770 233778
rect 589150 198098 589182 198334
rect 589418 198098 589502 198334
rect 589738 198098 589770 198334
rect 589150 198014 589770 198098
rect 589150 197778 589182 198014
rect 589418 197778 589502 198014
rect 589738 197778 589770 198014
rect 589150 162334 589770 197778
rect 589150 162098 589182 162334
rect 589418 162098 589502 162334
rect 589738 162098 589770 162334
rect 589150 162014 589770 162098
rect 589150 161778 589182 162014
rect 589418 161778 589502 162014
rect 589738 161778 589770 162014
rect 589150 126334 589770 161778
rect 589150 126098 589182 126334
rect 589418 126098 589502 126334
rect 589738 126098 589770 126334
rect 589150 126014 589770 126098
rect 589150 125778 589182 126014
rect 589418 125778 589502 126014
rect 589738 125778 589770 126014
rect 589150 90334 589770 125778
rect 589150 90098 589182 90334
rect 589418 90098 589502 90334
rect 589738 90098 589770 90334
rect 589150 90014 589770 90098
rect 589150 89778 589182 90014
rect 589418 89778 589502 90014
rect 589738 89778 589770 90014
rect 589150 54334 589770 89778
rect 589150 54098 589182 54334
rect 589418 54098 589502 54334
rect 589738 54098 589770 54334
rect 589150 54014 589770 54098
rect 589150 53778 589182 54014
rect 589418 53778 589502 54014
rect 589738 53778 589770 54014
rect 589150 18334 589770 53778
rect 589150 18098 589182 18334
rect 589418 18098 589502 18334
rect 589738 18098 589770 18334
rect 589150 18014 589770 18098
rect 589150 17778 589182 18014
rect 589418 17778 589502 18014
rect 589738 17778 589770 18014
rect 589150 -4186 589770 17778
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 670054 590730 709082
rect 590110 669818 590142 670054
rect 590378 669818 590462 670054
rect 590698 669818 590730 670054
rect 590110 669734 590730 669818
rect 590110 669498 590142 669734
rect 590378 669498 590462 669734
rect 590698 669498 590730 669734
rect 590110 634054 590730 669498
rect 590110 633818 590142 634054
rect 590378 633818 590462 634054
rect 590698 633818 590730 634054
rect 590110 633734 590730 633818
rect 590110 633498 590142 633734
rect 590378 633498 590462 633734
rect 590698 633498 590730 633734
rect 590110 598054 590730 633498
rect 590110 597818 590142 598054
rect 590378 597818 590462 598054
rect 590698 597818 590730 598054
rect 590110 597734 590730 597818
rect 590110 597498 590142 597734
rect 590378 597498 590462 597734
rect 590698 597498 590730 597734
rect 590110 562054 590730 597498
rect 590110 561818 590142 562054
rect 590378 561818 590462 562054
rect 590698 561818 590730 562054
rect 590110 561734 590730 561818
rect 590110 561498 590142 561734
rect 590378 561498 590462 561734
rect 590698 561498 590730 561734
rect 590110 526054 590730 561498
rect 590110 525818 590142 526054
rect 590378 525818 590462 526054
rect 590698 525818 590730 526054
rect 590110 525734 590730 525818
rect 590110 525498 590142 525734
rect 590378 525498 590462 525734
rect 590698 525498 590730 525734
rect 590110 490054 590730 525498
rect 590110 489818 590142 490054
rect 590378 489818 590462 490054
rect 590698 489818 590730 490054
rect 590110 489734 590730 489818
rect 590110 489498 590142 489734
rect 590378 489498 590462 489734
rect 590698 489498 590730 489734
rect 590110 454054 590730 489498
rect 590110 453818 590142 454054
rect 590378 453818 590462 454054
rect 590698 453818 590730 454054
rect 590110 453734 590730 453818
rect 590110 453498 590142 453734
rect 590378 453498 590462 453734
rect 590698 453498 590730 453734
rect 590110 418054 590730 453498
rect 590110 417818 590142 418054
rect 590378 417818 590462 418054
rect 590698 417818 590730 418054
rect 590110 417734 590730 417818
rect 590110 417498 590142 417734
rect 590378 417498 590462 417734
rect 590698 417498 590730 417734
rect 590110 382054 590730 417498
rect 590110 381818 590142 382054
rect 590378 381818 590462 382054
rect 590698 381818 590730 382054
rect 590110 381734 590730 381818
rect 590110 381498 590142 381734
rect 590378 381498 590462 381734
rect 590698 381498 590730 381734
rect 590110 346054 590730 381498
rect 590110 345818 590142 346054
rect 590378 345818 590462 346054
rect 590698 345818 590730 346054
rect 590110 345734 590730 345818
rect 590110 345498 590142 345734
rect 590378 345498 590462 345734
rect 590698 345498 590730 345734
rect 590110 310054 590730 345498
rect 590110 309818 590142 310054
rect 590378 309818 590462 310054
rect 590698 309818 590730 310054
rect 590110 309734 590730 309818
rect 590110 309498 590142 309734
rect 590378 309498 590462 309734
rect 590698 309498 590730 309734
rect 590110 274054 590730 309498
rect 590110 273818 590142 274054
rect 590378 273818 590462 274054
rect 590698 273818 590730 274054
rect 590110 273734 590730 273818
rect 590110 273498 590142 273734
rect 590378 273498 590462 273734
rect 590698 273498 590730 273734
rect 590110 238054 590730 273498
rect 590110 237818 590142 238054
rect 590378 237818 590462 238054
rect 590698 237818 590730 238054
rect 590110 237734 590730 237818
rect 590110 237498 590142 237734
rect 590378 237498 590462 237734
rect 590698 237498 590730 237734
rect 590110 202054 590730 237498
rect 590110 201818 590142 202054
rect 590378 201818 590462 202054
rect 590698 201818 590730 202054
rect 590110 201734 590730 201818
rect 590110 201498 590142 201734
rect 590378 201498 590462 201734
rect 590698 201498 590730 201734
rect 590110 166054 590730 201498
rect 590110 165818 590142 166054
rect 590378 165818 590462 166054
rect 590698 165818 590730 166054
rect 590110 165734 590730 165818
rect 590110 165498 590142 165734
rect 590378 165498 590462 165734
rect 590698 165498 590730 165734
rect 590110 130054 590730 165498
rect 590110 129818 590142 130054
rect 590378 129818 590462 130054
rect 590698 129818 590730 130054
rect 590110 129734 590730 129818
rect 590110 129498 590142 129734
rect 590378 129498 590462 129734
rect 590698 129498 590730 129734
rect 590110 94054 590730 129498
rect 590110 93818 590142 94054
rect 590378 93818 590462 94054
rect 590698 93818 590730 94054
rect 590110 93734 590730 93818
rect 590110 93498 590142 93734
rect 590378 93498 590462 93734
rect 590698 93498 590730 93734
rect 590110 58054 590730 93498
rect 590110 57818 590142 58054
rect 590378 57818 590462 58054
rect 590698 57818 590730 58054
rect 590110 57734 590730 57818
rect 590110 57498 590142 57734
rect 590378 57498 590462 57734
rect 590698 57498 590730 57734
rect 590110 22054 590730 57498
rect 590110 21818 590142 22054
rect 590378 21818 590462 22054
rect 590698 21818 590730 22054
rect 590110 21734 590730 21818
rect 590110 21498 590142 21734
rect 590378 21498 590462 21734
rect 590698 21498 590730 21734
rect 590110 -5146 590730 21498
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 673774 591690 710042
rect 591070 673538 591102 673774
rect 591338 673538 591422 673774
rect 591658 673538 591690 673774
rect 591070 673454 591690 673538
rect 591070 673218 591102 673454
rect 591338 673218 591422 673454
rect 591658 673218 591690 673454
rect 591070 637774 591690 673218
rect 591070 637538 591102 637774
rect 591338 637538 591422 637774
rect 591658 637538 591690 637774
rect 591070 637454 591690 637538
rect 591070 637218 591102 637454
rect 591338 637218 591422 637454
rect 591658 637218 591690 637454
rect 591070 601774 591690 637218
rect 591070 601538 591102 601774
rect 591338 601538 591422 601774
rect 591658 601538 591690 601774
rect 591070 601454 591690 601538
rect 591070 601218 591102 601454
rect 591338 601218 591422 601454
rect 591658 601218 591690 601454
rect 591070 565774 591690 601218
rect 591070 565538 591102 565774
rect 591338 565538 591422 565774
rect 591658 565538 591690 565774
rect 591070 565454 591690 565538
rect 591070 565218 591102 565454
rect 591338 565218 591422 565454
rect 591658 565218 591690 565454
rect 591070 529774 591690 565218
rect 591070 529538 591102 529774
rect 591338 529538 591422 529774
rect 591658 529538 591690 529774
rect 591070 529454 591690 529538
rect 591070 529218 591102 529454
rect 591338 529218 591422 529454
rect 591658 529218 591690 529454
rect 591070 493774 591690 529218
rect 591070 493538 591102 493774
rect 591338 493538 591422 493774
rect 591658 493538 591690 493774
rect 591070 493454 591690 493538
rect 591070 493218 591102 493454
rect 591338 493218 591422 493454
rect 591658 493218 591690 493454
rect 591070 457774 591690 493218
rect 591070 457538 591102 457774
rect 591338 457538 591422 457774
rect 591658 457538 591690 457774
rect 591070 457454 591690 457538
rect 591070 457218 591102 457454
rect 591338 457218 591422 457454
rect 591658 457218 591690 457454
rect 591070 421774 591690 457218
rect 591070 421538 591102 421774
rect 591338 421538 591422 421774
rect 591658 421538 591690 421774
rect 591070 421454 591690 421538
rect 591070 421218 591102 421454
rect 591338 421218 591422 421454
rect 591658 421218 591690 421454
rect 591070 385774 591690 421218
rect 591070 385538 591102 385774
rect 591338 385538 591422 385774
rect 591658 385538 591690 385774
rect 591070 385454 591690 385538
rect 591070 385218 591102 385454
rect 591338 385218 591422 385454
rect 591658 385218 591690 385454
rect 591070 349774 591690 385218
rect 591070 349538 591102 349774
rect 591338 349538 591422 349774
rect 591658 349538 591690 349774
rect 591070 349454 591690 349538
rect 591070 349218 591102 349454
rect 591338 349218 591422 349454
rect 591658 349218 591690 349454
rect 591070 313774 591690 349218
rect 591070 313538 591102 313774
rect 591338 313538 591422 313774
rect 591658 313538 591690 313774
rect 591070 313454 591690 313538
rect 591070 313218 591102 313454
rect 591338 313218 591422 313454
rect 591658 313218 591690 313454
rect 591070 277774 591690 313218
rect 591070 277538 591102 277774
rect 591338 277538 591422 277774
rect 591658 277538 591690 277774
rect 591070 277454 591690 277538
rect 591070 277218 591102 277454
rect 591338 277218 591422 277454
rect 591658 277218 591690 277454
rect 591070 241774 591690 277218
rect 591070 241538 591102 241774
rect 591338 241538 591422 241774
rect 591658 241538 591690 241774
rect 591070 241454 591690 241538
rect 591070 241218 591102 241454
rect 591338 241218 591422 241454
rect 591658 241218 591690 241454
rect 591070 205774 591690 241218
rect 591070 205538 591102 205774
rect 591338 205538 591422 205774
rect 591658 205538 591690 205774
rect 591070 205454 591690 205538
rect 591070 205218 591102 205454
rect 591338 205218 591422 205454
rect 591658 205218 591690 205454
rect 591070 169774 591690 205218
rect 591070 169538 591102 169774
rect 591338 169538 591422 169774
rect 591658 169538 591690 169774
rect 591070 169454 591690 169538
rect 591070 169218 591102 169454
rect 591338 169218 591422 169454
rect 591658 169218 591690 169454
rect 591070 133774 591690 169218
rect 591070 133538 591102 133774
rect 591338 133538 591422 133774
rect 591658 133538 591690 133774
rect 591070 133454 591690 133538
rect 591070 133218 591102 133454
rect 591338 133218 591422 133454
rect 591658 133218 591690 133454
rect 591070 97774 591690 133218
rect 591070 97538 591102 97774
rect 591338 97538 591422 97774
rect 591658 97538 591690 97774
rect 591070 97454 591690 97538
rect 591070 97218 591102 97454
rect 591338 97218 591422 97454
rect 591658 97218 591690 97454
rect 591070 61774 591690 97218
rect 591070 61538 591102 61774
rect 591338 61538 591422 61774
rect 591658 61538 591690 61774
rect 591070 61454 591690 61538
rect 591070 61218 591102 61454
rect 591338 61218 591422 61454
rect 591658 61218 591690 61454
rect 591070 25774 591690 61218
rect 591070 25538 591102 25774
rect 591338 25538 591422 25774
rect 591658 25538 591690 25774
rect 591070 25454 591690 25538
rect 591070 25218 591102 25454
rect 591338 25218 591422 25454
rect 591658 25218 591690 25454
rect 591070 -6106 591690 25218
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 677494 592650 711002
rect 592030 677258 592062 677494
rect 592298 677258 592382 677494
rect 592618 677258 592650 677494
rect 592030 677174 592650 677258
rect 592030 676938 592062 677174
rect 592298 676938 592382 677174
rect 592618 676938 592650 677174
rect 592030 641494 592650 676938
rect 592030 641258 592062 641494
rect 592298 641258 592382 641494
rect 592618 641258 592650 641494
rect 592030 641174 592650 641258
rect 592030 640938 592062 641174
rect 592298 640938 592382 641174
rect 592618 640938 592650 641174
rect 592030 605494 592650 640938
rect 592030 605258 592062 605494
rect 592298 605258 592382 605494
rect 592618 605258 592650 605494
rect 592030 605174 592650 605258
rect 592030 604938 592062 605174
rect 592298 604938 592382 605174
rect 592618 604938 592650 605174
rect 592030 569494 592650 604938
rect 592030 569258 592062 569494
rect 592298 569258 592382 569494
rect 592618 569258 592650 569494
rect 592030 569174 592650 569258
rect 592030 568938 592062 569174
rect 592298 568938 592382 569174
rect 592618 568938 592650 569174
rect 592030 533494 592650 568938
rect 592030 533258 592062 533494
rect 592298 533258 592382 533494
rect 592618 533258 592650 533494
rect 592030 533174 592650 533258
rect 592030 532938 592062 533174
rect 592298 532938 592382 533174
rect 592618 532938 592650 533174
rect 592030 497494 592650 532938
rect 592030 497258 592062 497494
rect 592298 497258 592382 497494
rect 592618 497258 592650 497494
rect 592030 497174 592650 497258
rect 592030 496938 592062 497174
rect 592298 496938 592382 497174
rect 592618 496938 592650 497174
rect 592030 461494 592650 496938
rect 592030 461258 592062 461494
rect 592298 461258 592382 461494
rect 592618 461258 592650 461494
rect 592030 461174 592650 461258
rect 592030 460938 592062 461174
rect 592298 460938 592382 461174
rect 592618 460938 592650 461174
rect 592030 425494 592650 460938
rect 592030 425258 592062 425494
rect 592298 425258 592382 425494
rect 592618 425258 592650 425494
rect 592030 425174 592650 425258
rect 592030 424938 592062 425174
rect 592298 424938 592382 425174
rect 592618 424938 592650 425174
rect 592030 389494 592650 424938
rect 592030 389258 592062 389494
rect 592298 389258 592382 389494
rect 592618 389258 592650 389494
rect 592030 389174 592650 389258
rect 592030 388938 592062 389174
rect 592298 388938 592382 389174
rect 592618 388938 592650 389174
rect 592030 353494 592650 388938
rect 592030 353258 592062 353494
rect 592298 353258 592382 353494
rect 592618 353258 592650 353494
rect 592030 353174 592650 353258
rect 592030 352938 592062 353174
rect 592298 352938 592382 353174
rect 592618 352938 592650 353174
rect 592030 317494 592650 352938
rect 592030 317258 592062 317494
rect 592298 317258 592382 317494
rect 592618 317258 592650 317494
rect 592030 317174 592650 317258
rect 592030 316938 592062 317174
rect 592298 316938 592382 317174
rect 592618 316938 592650 317174
rect 592030 281494 592650 316938
rect 592030 281258 592062 281494
rect 592298 281258 592382 281494
rect 592618 281258 592650 281494
rect 592030 281174 592650 281258
rect 592030 280938 592062 281174
rect 592298 280938 592382 281174
rect 592618 280938 592650 281174
rect 592030 245494 592650 280938
rect 592030 245258 592062 245494
rect 592298 245258 592382 245494
rect 592618 245258 592650 245494
rect 592030 245174 592650 245258
rect 592030 244938 592062 245174
rect 592298 244938 592382 245174
rect 592618 244938 592650 245174
rect 592030 209494 592650 244938
rect 592030 209258 592062 209494
rect 592298 209258 592382 209494
rect 592618 209258 592650 209494
rect 592030 209174 592650 209258
rect 592030 208938 592062 209174
rect 592298 208938 592382 209174
rect 592618 208938 592650 209174
rect 592030 173494 592650 208938
rect 592030 173258 592062 173494
rect 592298 173258 592382 173494
rect 592618 173258 592650 173494
rect 592030 173174 592650 173258
rect 592030 172938 592062 173174
rect 592298 172938 592382 173174
rect 592618 172938 592650 173174
rect 592030 137494 592650 172938
rect 592030 137258 592062 137494
rect 592298 137258 592382 137494
rect 592618 137258 592650 137494
rect 592030 137174 592650 137258
rect 592030 136938 592062 137174
rect 592298 136938 592382 137174
rect 592618 136938 592650 137174
rect 592030 101494 592650 136938
rect 592030 101258 592062 101494
rect 592298 101258 592382 101494
rect 592618 101258 592650 101494
rect 592030 101174 592650 101258
rect 592030 100938 592062 101174
rect 592298 100938 592382 101174
rect 592618 100938 592650 101174
rect 592030 65494 592650 100938
rect 592030 65258 592062 65494
rect 592298 65258 592382 65494
rect 592618 65258 592650 65494
rect 592030 65174 592650 65258
rect 592030 64938 592062 65174
rect 592298 64938 592382 65174
rect 592618 64938 592650 65174
rect 592030 29494 592650 64938
rect 592030 29258 592062 29494
rect 592298 29258 592382 29494
rect 592618 29258 592650 29494
rect 592030 29174 592650 29258
rect 592030 28938 592062 29174
rect 592298 28938 592382 29174
rect 592618 28938 592650 29174
rect 592030 -7066 592650 28938
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 677258 -8458 677494
rect -8374 677258 -8138 677494
rect -8694 676938 -8458 677174
rect -8374 676938 -8138 677174
rect -8694 641258 -8458 641494
rect -8374 641258 -8138 641494
rect -8694 640938 -8458 641174
rect -8374 640938 -8138 641174
rect -8694 605258 -8458 605494
rect -8374 605258 -8138 605494
rect -8694 604938 -8458 605174
rect -8374 604938 -8138 605174
rect -8694 569258 -8458 569494
rect -8374 569258 -8138 569494
rect -8694 568938 -8458 569174
rect -8374 568938 -8138 569174
rect -8694 533258 -8458 533494
rect -8374 533258 -8138 533494
rect -8694 532938 -8458 533174
rect -8374 532938 -8138 533174
rect -8694 497258 -8458 497494
rect -8374 497258 -8138 497494
rect -8694 496938 -8458 497174
rect -8374 496938 -8138 497174
rect -8694 461258 -8458 461494
rect -8374 461258 -8138 461494
rect -8694 460938 -8458 461174
rect -8374 460938 -8138 461174
rect -8694 425258 -8458 425494
rect -8374 425258 -8138 425494
rect -8694 424938 -8458 425174
rect -8374 424938 -8138 425174
rect -8694 389258 -8458 389494
rect -8374 389258 -8138 389494
rect -8694 388938 -8458 389174
rect -8374 388938 -8138 389174
rect -8694 353258 -8458 353494
rect -8374 353258 -8138 353494
rect -8694 352938 -8458 353174
rect -8374 352938 -8138 353174
rect -8694 317258 -8458 317494
rect -8374 317258 -8138 317494
rect -8694 316938 -8458 317174
rect -8374 316938 -8138 317174
rect -8694 281258 -8458 281494
rect -8374 281258 -8138 281494
rect -8694 280938 -8458 281174
rect -8374 280938 -8138 281174
rect -8694 245258 -8458 245494
rect -8374 245258 -8138 245494
rect -8694 244938 -8458 245174
rect -8374 244938 -8138 245174
rect -8694 209258 -8458 209494
rect -8374 209258 -8138 209494
rect -8694 208938 -8458 209174
rect -8374 208938 -8138 209174
rect -8694 173258 -8458 173494
rect -8374 173258 -8138 173494
rect -8694 172938 -8458 173174
rect -8374 172938 -8138 173174
rect -8694 137258 -8458 137494
rect -8374 137258 -8138 137494
rect -8694 136938 -8458 137174
rect -8374 136938 -8138 137174
rect -8694 101258 -8458 101494
rect -8374 101258 -8138 101494
rect -8694 100938 -8458 101174
rect -8374 100938 -8138 101174
rect -8694 65258 -8458 65494
rect -8374 65258 -8138 65494
rect -8694 64938 -8458 65174
rect -8374 64938 -8138 65174
rect -8694 29258 -8458 29494
rect -8374 29258 -8138 29494
rect -8694 28938 -8458 29174
rect -8374 28938 -8138 29174
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 673538 -7498 673774
rect -7414 673538 -7178 673774
rect -7734 673218 -7498 673454
rect -7414 673218 -7178 673454
rect -7734 637538 -7498 637774
rect -7414 637538 -7178 637774
rect -7734 637218 -7498 637454
rect -7414 637218 -7178 637454
rect -7734 601538 -7498 601774
rect -7414 601538 -7178 601774
rect -7734 601218 -7498 601454
rect -7414 601218 -7178 601454
rect -7734 565538 -7498 565774
rect -7414 565538 -7178 565774
rect -7734 565218 -7498 565454
rect -7414 565218 -7178 565454
rect -7734 529538 -7498 529774
rect -7414 529538 -7178 529774
rect -7734 529218 -7498 529454
rect -7414 529218 -7178 529454
rect -7734 493538 -7498 493774
rect -7414 493538 -7178 493774
rect -7734 493218 -7498 493454
rect -7414 493218 -7178 493454
rect -7734 457538 -7498 457774
rect -7414 457538 -7178 457774
rect -7734 457218 -7498 457454
rect -7414 457218 -7178 457454
rect -7734 421538 -7498 421774
rect -7414 421538 -7178 421774
rect -7734 421218 -7498 421454
rect -7414 421218 -7178 421454
rect -7734 385538 -7498 385774
rect -7414 385538 -7178 385774
rect -7734 385218 -7498 385454
rect -7414 385218 -7178 385454
rect -7734 349538 -7498 349774
rect -7414 349538 -7178 349774
rect -7734 349218 -7498 349454
rect -7414 349218 -7178 349454
rect -7734 313538 -7498 313774
rect -7414 313538 -7178 313774
rect -7734 313218 -7498 313454
rect -7414 313218 -7178 313454
rect -7734 277538 -7498 277774
rect -7414 277538 -7178 277774
rect -7734 277218 -7498 277454
rect -7414 277218 -7178 277454
rect -7734 241538 -7498 241774
rect -7414 241538 -7178 241774
rect -7734 241218 -7498 241454
rect -7414 241218 -7178 241454
rect -7734 205538 -7498 205774
rect -7414 205538 -7178 205774
rect -7734 205218 -7498 205454
rect -7414 205218 -7178 205454
rect -7734 169538 -7498 169774
rect -7414 169538 -7178 169774
rect -7734 169218 -7498 169454
rect -7414 169218 -7178 169454
rect -7734 133538 -7498 133774
rect -7414 133538 -7178 133774
rect -7734 133218 -7498 133454
rect -7414 133218 -7178 133454
rect -7734 97538 -7498 97774
rect -7414 97538 -7178 97774
rect -7734 97218 -7498 97454
rect -7414 97218 -7178 97454
rect -7734 61538 -7498 61774
rect -7414 61538 -7178 61774
rect -7734 61218 -7498 61454
rect -7414 61218 -7178 61454
rect -7734 25538 -7498 25774
rect -7414 25538 -7178 25774
rect -7734 25218 -7498 25454
rect -7414 25218 -7178 25454
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 669818 -6538 670054
rect -6454 669818 -6218 670054
rect -6774 669498 -6538 669734
rect -6454 669498 -6218 669734
rect -6774 633818 -6538 634054
rect -6454 633818 -6218 634054
rect -6774 633498 -6538 633734
rect -6454 633498 -6218 633734
rect -6774 597818 -6538 598054
rect -6454 597818 -6218 598054
rect -6774 597498 -6538 597734
rect -6454 597498 -6218 597734
rect -6774 561818 -6538 562054
rect -6454 561818 -6218 562054
rect -6774 561498 -6538 561734
rect -6454 561498 -6218 561734
rect -6774 525818 -6538 526054
rect -6454 525818 -6218 526054
rect -6774 525498 -6538 525734
rect -6454 525498 -6218 525734
rect -6774 489818 -6538 490054
rect -6454 489818 -6218 490054
rect -6774 489498 -6538 489734
rect -6454 489498 -6218 489734
rect -6774 453818 -6538 454054
rect -6454 453818 -6218 454054
rect -6774 453498 -6538 453734
rect -6454 453498 -6218 453734
rect -6774 417818 -6538 418054
rect -6454 417818 -6218 418054
rect -6774 417498 -6538 417734
rect -6454 417498 -6218 417734
rect -6774 381818 -6538 382054
rect -6454 381818 -6218 382054
rect -6774 381498 -6538 381734
rect -6454 381498 -6218 381734
rect -6774 345818 -6538 346054
rect -6454 345818 -6218 346054
rect -6774 345498 -6538 345734
rect -6454 345498 -6218 345734
rect -6774 309818 -6538 310054
rect -6454 309818 -6218 310054
rect -6774 309498 -6538 309734
rect -6454 309498 -6218 309734
rect -6774 273818 -6538 274054
rect -6454 273818 -6218 274054
rect -6774 273498 -6538 273734
rect -6454 273498 -6218 273734
rect -6774 237818 -6538 238054
rect -6454 237818 -6218 238054
rect -6774 237498 -6538 237734
rect -6454 237498 -6218 237734
rect -6774 201818 -6538 202054
rect -6454 201818 -6218 202054
rect -6774 201498 -6538 201734
rect -6454 201498 -6218 201734
rect -6774 165818 -6538 166054
rect -6454 165818 -6218 166054
rect -6774 165498 -6538 165734
rect -6454 165498 -6218 165734
rect -6774 129818 -6538 130054
rect -6454 129818 -6218 130054
rect -6774 129498 -6538 129734
rect -6454 129498 -6218 129734
rect -6774 93818 -6538 94054
rect -6454 93818 -6218 94054
rect -6774 93498 -6538 93734
rect -6454 93498 -6218 93734
rect -6774 57818 -6538 58054
rect -6454 57818 -6218 58054
rect -6774 57498 -6538 57734
rect -6454 57498 -6218 57734
rect -6774 21818 -6538 22054
rect -6454 21818 -6218 22054
rect -6774 21498 -6538 21734
rect -6454 21498 -6218 21734
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 666098 -5578 666334
rect -5494 666098 -5258 666334
rect -5814 665778 -5578 666014
rect -5494 665778 -5258 666014
rect -5814 630098 -5578 630334
rect -5494 630098 -5258 630334
rect -5814 629778 -5578 630014
rect -5494 629778 -5258 630014
rect -5814 594098 -5578 594334
rect -5494 594098 -5258 594334
rect -5814 593778 -5578 594014
rect -5494 593778 -5258 594014
rect -5814 558098 -5578 558334
rect -5494 558098 -5258 558334
rect -5814 557778 -5578 558014
rect -5494 557778 -5258 558014
rect -5814 522098 -5578 522334
rect -5494 522098 -5258 522334
rect -5814 521778 -5578 522014
rect -5494 521778 -5258 522014
rect -5814 486098 -5578 486334
rect -5494 486098 -5258 486334
rect -5814 485778 -5578 486014
rect -5494 485778 -5258 486014
rect -5814 450098 -5578 450334
rect -5494 450098 -5258 450334
rect -5814 449778 -5578 450014
rect -5494 449778 -5258 450014
rect -5814 414098 -5578 414334
rect -5494 414098 -5258 414334
rect -5814 413778 -5578 414014
rect -5494 413778 -5258 414014
rect -5814 378098 -5578 378334
rect -5494 378098 -5258 378334
rect -5814 377778 -5578 378014
rect -5494 377778 -5258 378014
rect -5814 342098 -5578 342334
rect -5494 342098 -5258 342334
rect -5814 341778 -5578 342014
rect -5494 341778 -5258 342014
rect -5814 306098 -5578 306334
rect -5494 306098 -5258 306334
rect -5814 305778 -5578 306014
rect -5494 305778 -5258 306014
rect -5814 270098 -5578 270334
rect -5494 270098 -5258 270334
rect -5814 269778 -5578 270014
rect -5494 269778 -5258 270014
rect -5814 234098 -5578 234334
rect -5494 234098 -5258 234334
rect -5814 233778 -5578 234014
rect -5494 233778 -5258 234014
rect -5814 198098 -5578 198334
rect -5494 198098 -5258 198334
rect -5814 197778 -5578 198014
rect -5494 197778 -5258 198014
rect -5814 162098 -5578 162334
rect -5494 162098 -5258 162334
rect -5814 161778 -5578 162014
rect -5494 161778 -5258 162014
rect -5814 126098 -5578 126334
rect -5494 126098 -5258 126334
rect -5814 125778 -5578 126014
rect -5494 125778 -5258 126014
rect -5814 90098 -5578 90334
rect -5494 90098 -5258 90334
rect -5814 89778 -5578 90014
rect -5494 89778 -5258 90014
rect -5814 54098 -5578 54334
rect -5494 54098 -5258 54334
rect -5814 53778 -5578 54014
rect -5494 53778 -5258 54014
rect -5814 18098 -5578 18334
rect -5494 18098 -5258 18334
rect -5814 17778 -5578 18014
rect -5494 17778 -5258 18014
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 698378 -4618 698614
rect -4534 698378 -4298 698614
rect -4854 698058 -4618 698294
rect -4534 698058 -4298 698294
rect -4854 662378 -4618 662614
rect -4534 662378 -4298 662614
rect -4854 662058 -4618 662294
rect -4534 662058 -4298 662294
rect -4854 626378 -4618 626614
rect -4534 626378 -4298 626614
rect -4854 626058 -4618 626294
rect -4534 626058 -4298 626294
rect -4854 590378 -4618 590614
rect -4534 590378 -4298 590614
rect -4854 590058 -4618 590294
rect -4534 590058 -4298 590294
rect -4854 554378 -4618 554614
rect -4534 554378 -4298 554614
rect -4854 554058 -4618 554294
rect -4534 554058 -4298 554294
rect -4854 518378 -4618 518614
rect -4534 518378 -4298 518614
rect -4854 518058 -4618 518294
rect -4534 518058 -4298 518294
rect -4854 482378 -4618 482614
rect -4534 482378 -4298 482614
rect -4854 482058 -4618 482294
rect -4534 482058 -4298 482294
rect -4854 446378 -4618 446614
rect -4534 446378 -4298 446614
rect -4854 446058 -4618 446294
rect -4534 446058 -4298 446294
rect -4854 410378 -4618 410614
rect -4534 410378 -4298 410614
rect -4854 410058 -4618 410294
rect -4534 410058 -4298 410294
rect -4854 374378 -4618 374614
rect -4534 374378 -4298 374614
rect -4854 374058 -4618 374294
rect -4534 374058 -4298 374294
rect -4854 338378 -4618 338614
rect -4534 338378 -4298 338614
rect -4854 338058 -4618 338294
rect -4534 338058 -4298 338294
rect -4854 302378 -4618 302614
rect -4534 302378 -4298 302614
rect -4854 302058 -4618 302294
rect -4534 302058 -4298 302294
rect -4854 266378 -4618 266614
rect -4534 266378 -4298 266614
rect -4854 266058 -4618 266294
rect -4534 266058 -4298 266294
rect -4854 230378 -4618 230614
rect -4534 230378 -4298 230614
rect -4854 230058 -4618 230294
rect -4534 230058 -4298 230294
rect -4854 194378 -4618 194614
rect -4534 194378 -4298 194614
rect -4854 194058 -4618 194294
rect -4534 194058 -4298 194294
rect -4854 158378 -4618 158614
rect -4534 158378 -4298 158614
rect -4854 158058 -4618 158294
rect -4534 158058 -4298 158294
rect -4854 122378 -4618 122614
rect -4534 122378 -4298 122614
rect -4854 122058 -4618 122294
rect -4534 122058 -4298 122294
rect -4854 86378 -4618 86614
rect -4534 86378 -4298 86614
rect -4854 86058 -4618 86294
rect -4534 86058 -4298 86294
rect -4854 50378 -4618 50614
rect -4534 50378 -4298 50614
rect -4854 50058 -4618 50294
rect -4534 50058 -4298 50294
rect -4854 14378 -4618 14614
rect -4534 14378 -4298 14614
rect -4854 14058 -4618 14294
rect -4534 14058 -4298 14294
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 694658 -3658 694894
rect -3574 694658 -3338 694894
rect -3894 694338 -3658 694574
rect -3574 694338 -3338 694574
rect -3894 658658 -3658 658894
rect -3574 658658 -3338 658894
rect -3894 658338 -3658 658574
rect -3574 658338 -3338 658574
rect -3894 622658 -3658 622894
rect -3574 622658 -3338 622894
rect -3894 622338 -3658 622574
rect -3574 622338 -3338 622574
rect -3894 586658 -3658 586894
rect -3574 586658 -3338 586894
rect -3894 586338 -3658 586574
rect -3574 586338 -3338 586574
rect -3894 550658 -3658 550894
rect -3574 550658 -3338 550894
rect -3894 550338 -3658 550574
rect -3574 550338 -3338 550574
rect -3894 514658 -3658 514894
rect -3574 514658 -3338 514894
rect -3894 514338 -3658 514574
rect -3574 514338 -3338 514574
rect -3894 478658 -3658 478894
rect -3574 478658 -3338 478894
rect -3894 478338 -3658 478574
rect -3574 478338 -3338 478574
rect -3894 442658 -3658 442894
rect -3574 442658 -3338 442894
rect -3894 442338 -3658 442574
rect -3574 442338 -3338 442574
rect -3894 406658 -3658 406894
rect -3574 406658 -3338 406894
rect -3894 406338 -3658 406574
rect -3574 406338 -3338 406574
rect -3894 370658 -3658 370894
rect -3574 370658 -3338 370894
rect -3894 370338 -3658 370574
rect -3574 370338 -3338 370574
rect -3894 334658 -3658 334894
rect -3574 334658 -3338 334894
rect -3894 334338 -3658 334574
rect -3574 334338 -3338 334574
rect -3894 298658 -3658 298894
rect -3574 298658 -3338 298894
rect -3894 298338 -3658 298574
rect -3574 298338 -3338 298574
rect -3894 262658 -3658 262894
rect -3574 262658 -3338 262894
rect -3894 262338 -3658 262574
rect -3574 262338 -3338 262574
rect -3894 226658 -3658 226894
rect -3574 226658 -3338 226894
rect -3894 226338 -3658 226574
rect -3574 226338 -3338 226574
rect -3894 190658 -3658 190894
rect -3574 190658 -3338 190894
rect -3894 190338 -3658 190574
rect -3574 190338 -3338 190574
rect -3894 154658 -3658 154894
rect -3574 154658 -3338 154894
rect -3894 154338 -3658 154574
rect -3574 154338 -3338 154574
rect -3894 118658 -3658 118894
rect -3574 118658 -3338 118894
rect -3894 118338 -3658 118574
rect -3574 118338 -3338 118574
rect -3894 82658 -3658 82894
rect -3574 82658 -3338 82894
rect -3894 82338 -3658 82574
rect -3574 82338 -3338 82574
rect -3894 46658 -3658 46894
rect -3574 46658 -3338 46894
rect -3894 46338 -3658 46574
rect -3574 46338 -3338 46574
rect -3894 10658 -3658 10894
rect -3574 10658 -3338 10894
rect -3894 10338 -3658 10574
rect -3574 10338 -3338 10574
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 690938 -2698 691174
rect -2614 690938 -2378 691174
rect -2934 690618 -2698 690854
rect -2614 690618 -2378 690854
rect -2934 654938 -2698 655174
rect -2614 654938 -2378 655174
rect -2934 654618 -2698 654854
rect -2614 654618 -2378 654854
rect -2934 618938 -2698 619174
rect -2614 618938 -2378 619174
rect -2934 618618 -2698 618854
rect -2614 618618 -2378 618854
rect -2934 582938 -2698 583174
rect -2614 582938 -2378 583174
rect -2934 582618 -2698 582854
rect -2614 582618 -2378 582854
rect -2934 546938 -2698 547174
rect -2614 546938 -2378 547174
rect -2934 546618 -2698 546854
rect -2614 546618 -2378 546854
rect -2934 510938 -2698 511174
rect -2614 510938 -2378 511174
rect -2934 510618 -2698 510854
rect -2614 510618 -2378 510854
rect -2934 474938 -2698 475174
rect -2614 474938 -2378 475174
rect -2934 474618 -2698 474854
rect -2614 474618 -2378 474854
rect -2934 438938 -2698 439174
rect -2614 438938 -2378 439174
rect -2934 438618 -2698 438854
rect -2614 438618 -2378 438854
rect -2934 402938 -2698 403174
rect -2614 402938 -2378 403174
rect -2934 402618 -2698 402854
rect -2614 402618 -2378 402854
rect -2934 366938 -2698 367174
rect -2614 366938 -2378 367174
rect -2934 366618 -2698 366854
rect -2614 366618 -2378 366854
rect -2934 330938 -2698 331174
rect -2614 330938 -2378 331174
rect -2934 330618 -2698 330854
rect -2614 330618 -2378 330854
rect -2934 294938 -2698 295174
rect -2614 294938 -2378 295174
rect -2934 294618 -2698 294854
rect -2614 294618 -2378 294854
rect -2934 258938 -2698 259174
rect -2614 258938 -2378 259174
rect -2934 258618 -2698 258854
rect -2614 258618 -2378 258854
rect -2934 222938 -2698 223174
rect -2614 222938 -2378 223174
rect -2934 222618 -2698 222854
rect -2614 222618 -2378 222854
rect -2934 186938 -2698 187174
rect -2614 186938 -2378 187174
rect -2934 186618 -2698 186854
rect -2614 186618 -2378 186854
rect -2934 150938 -2698 151174
rect -2614 150938 -2378 151174
rect -2934 150618 -2698 150854
rect -2614 150618 -2378 150854
rect -2934 114938 -2698 115174
rect -2614 114938 -2378 115174
rect -2934 114618 -2698 114854
rect -2614 114618 -2378 114854
rect -2934 78938 -2698 79174
rect -2614 78938 -2378 79174
rect -2934 78618 -2698 78854
rect -2614 78618 -2378 78854
rect -2934 42938 -2698 43174
rect -2614 42938 -2378 43174
rect -2934 42618 -2698 42854
rect -2614 42618 -2378 42854
rect -2934 6938 -2698 7174
rect -2614 6938 -2378 7174
rect -2934 6618 -2698 6854
rect -2614 6618 -2378 6854
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 9266 706522 9502 706758
rect 9586 706522 9822 706758
rect 9266 706202 9502 706438
rect 9586 706202 9822 706438
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 12986 707482 13222 707718
rect 13306 707482 13542 707718
rect 12986 707162 13222 707398
rect 13306 707162 13542 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 45266 706522 45502 706758
rect 45586 706522 45822 706758
rect 45266 706202 45502 706438
rect 45586 706202 45822 706438
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 48986 707482 49222 707718
rect 49306 707482 49542 707718
rect 48986 707162 49222 707398
rect 49306 707162 49542 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 81266 706522 81502 706758
rect 81586 706522 81822 706758
rect 81266 706202 81502 706438
rect 81586 706202 81822 706438
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 84986 707482 85222 707718
rect 85306 707482 85542 707718
rect 84986 707162 85222 707398
rect 85306 707162 85542 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 117266 706522 117502 706758
rect 117586 706522 117822 706758
rect 117266 706202 117502 706438
rect 117586 706202 117822 706438
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 120986 707482 121222 707718
rect 121306 707482 121542 707718
rect 120986 707162 121222 707398
rect 121306 707162 121542 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 153266 706522 153502 706758
rect 153586 706522 153822 706758
rect 153266 706202 153502 706438
rect 153586 706202 153822 706438
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 156986 707482 157222 707718
rect 157306 707482 157542 707718
rect 156986 707162 157222 707398
rect 157306 707162 157542 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 189266 706522 189502 706758
rect 189586 706522 189822 706758
rect 189266 706202 189502 706438
rect 189586 706202 189822 706438
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 192986 707482 193222 707718
rect 193306 707482 193542 707718
rect 192986 707162 193222 707398
rect 193306 707162 193542 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 225266 706522 225502 706758
rect 225586 706522 225822 706758
rect 225266 706202 225502 706438
rect 225586 706202 225822 706438
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 228986 707482 229222 707718
rect 229306 707482 229542 707718
rect 228986 707162 229222 707398
rect 229306 707162 229542 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 261266 706522 261502 706758
rect 261586 706522 261822 706758
rect 261266 706202 261502 706438
rect 261586 706202 261822 706438
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 264986 707482 265222 707718
rect 265306 707482 265542 707718
rect 264986 707162 265222 707398
rect 265306 707162 265542 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 297266 706522 297502 706758
rect 297586 706522 297822 706758
rect 297266 706202 297502 706438
rect 297586 706202 297822 706438
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 300986 707482 301222 707718
rect 301306 707482 301542 707718
rect 300986 707162 301222 707398
rect 301306 707162 301542 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 333266 706522 333502 706758
rect 333586 706522 333822 706758
rect 333266 706202 333502 706438
rect 333586 706202 333822 706438
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 336986 707482 337222 707718
rect 337306 707482 337542 707718
rect 336986 707162 337222 707398
rect 337306 707162 337542 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 369266 706522 369502 706758
rect 369586 706522 369822 706758
rect 369266 706202 369502 706438
rect 369586 706202 369822 706438
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 372986 707482 373222 707718
rect 373306 707482 373542 707718
rect 372986 707162 373222 707398
rect 373306 707162 373542 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 405266 706522 405502 706758
rect 405586 706522 405822 706758
rect 405266 706202 405502 706438
rect 405586 706202 405822 706438
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 408986 707482 409222 707718
rect 409306 707482 409542 707718
rect 408986 707162 409222 707398
rect 409306 707162 409542 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 441266 706522 441502 706758
rect 441586 706522 441822 706758
rect 441266 706202 441502 706438
rect 441586 706202 441822 706438
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 444986 707482 445222 707718
rect 445306 707482 445542 707718
rect 444986 707162 445222 707398
rect 445306 707162 445542 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 477266 706522 477502 706758
rect 477586 706522 477822 706758
rect 477266 706202 477502 706438
rect 477586 706202 477822 706438
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 480986 707482 481222 707718
rect 481306 707482 481542 707718
rect 480986 707162 481222 707398
rect 481306 707162 481542 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 513266 706522 513502 706758
rect 513586 706522 513822 706758
rect 513266 706202 513502 706438
rect 513586 706202 513822 706438
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 516986 707482 517222 707718
rect 517306 707482 517542 707718
rect 516986 707162 517222 707398
rect 517306 707162 517542 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 549266 706522 549502 706758
rect 549586 706522 549822 706758
rect 549266 706202 549502 706438
rect 549586 706202 549822 706438
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 552986 707482 553222 707718
rect 553306 707482 553542 707718
rect 552986 707162 553222 707398
rect 553306 707162 553542 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 10250 687218 10486 687454
rect 10250 686898 10486 687134
rect 40970 687218 41206 687454
rect 40970 686898 41206 687134
rect 71690 687218 71926 687454
rect 71690 686898 71926 687134
rect 102410 687218 102646 687454
rect 102410 686898 102646 687134
rect 133130 687218 133366 687454
rect 133130 686898 133366 687134
rect 163850 687218 164086 687454
rect 163850 686898 164086 687134
rect 194570 687218 194806 687454
rect 194570 686898 194806 687134
rect 225290 687218 225526 687454
rect 225290 686898 225526 687134
rect 256010 687218 256246 687454
rect 256010 686898 256246 687134
rect 286730 687218 286966 687454
rect 286730 686898 286966 687134
rect 317450 687218 317686 687454
rect 317450 686898 317686 687134
rect 348170 687218 348406 687454
rect 348170 686898 348406 687134
rect 378890 687218 379126 687454
rect 378890 686898 379126 687134
rect 409610 687218 409846 687454
rect 409610 686898 409846 687134
rect 440330 687218 440566 687454
rect 440330 686898 440566 687134
rect 471050 687218 471286 687454
rect 471050 686898 471286 687134
rect 501770 687218 502006 687454
rect 501770 686898 502006 687134
rect 532490 687218 532726 687454
rect 532490 686898 532726 687134
rect 563210 687218 563446 687454
rect 563210 686898 563446 687134
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 25610 654938 25846 655174
rect 25610 654618 25846 654854
rect 56330 654938 56566 655174
rect 56330 654618 56566 654854
rect 87050 654938 87286 655174
rect 87050 654618 87286 654854
rect 117770 654938 118006 655174
rect 117770 654618 118006 654854
rect 148490 654938 148726 655174
rect 148490 654618 148726 654854
rect 179210 654938 179446 655174
rect 179210 654618 179446 654854
rect 209930 654938 210166 655174
rect 209930 654618 210166 654854
rect 240650 654938 240886 655174
rect 240650 654618 240886 654854
rect 271370 654938 271606 655174
rect 271370 654618 271606 654854
rect 302090 654938 302326 655174
rect 302090 654618 302326 654854
rect 332810 654938 333046 655174
rect 332810 654618 333046 654854
rect 363530 654938 363766 655174
rect 363530 654618 363766 654854
rect 394250 654938 394486 655174
rect 394250 654618 394486 654854
rect 424970 654938 425206 655174
rect 424970 654618 425206 654854
rect 455690 654938 455926 655174
rect 455690 654618 455926 654854
rect 486410 654938 486646 655174
rect 486410 654618 486646 654854
rect 517130 654938 517366 655174
rect 517130 654618 517366 654854
rect 547850 654938 548086 655174
rect 547850 654618 548086 654854
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 10250 651218 10486 651454
rect 10250 650898 10486 651134
rect 40970 651218 41206 651454
rect 40970 650898 41206 651134
rect 71690 651218 71926 651454
rect 71690 650898 71926 651134
rect 102410 651218 102646 651454
rect 102410 650898 102646 651134
rect 133130 651218 133366 651454
rect 133130 650898 133366 651134
rect 163850 651218 164086 651454
rect 163850 650898 164086 651134
rect 194570 651218 194806 651454
rect 194570 650898 194806 651134
rect 225290 651218 225526 651454
rect 225290 650898 225526 651134
rect 256010 651218 256246 651454
rect 256010 650898 256246 651134
rect 286730 651218 286966 651454
rect 286730 650898 286966 651134
rect 317450 651218 317686 651454
rect 317450 650898 317686 651134
rect 348170 651218 348406 651454
rect 348170 650898 348406 651134
rect 378890 651218 379126 651454
rect 378890 650898 379126 651134
rect 409610 651218 409846 651454
rect 409610 650898 409846 651134
rect 440330 651218 440566 651454
rect 440330 650898 440566 651134
rect 471050 651218 471286 651454
rect 471050 650898 471286 651134
rect 501770 651218 502006 651454
rect 501770 650898 502006 651134
rect 532490 651218 532726 651454
rect 532490 650898 532726 651134
rect 563210 651218 563446 651454
rect 563210 650898 563446 651134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 25610 618938 25846 619174
rect 25610 618618 25846 618854
rect 56330 618938 56566 619174
rect 56330 618618 56566 618854
rect 87050 618938 87286 619174
rect 87050 618618 87286 618854
rect 117770 618938 118006 619174
rect 117770 618618 118006 618854
rect 148490 618938 148726 619174
rect 148490 618618 148726 618854
rect 179210 618938 179446 619174
rect 179210 618618 179446 618854
rect 209930 618938 210166 619174
rect 209930 618618 210166 618854
rect 240650 618938 240886 619174
rect 240650 618618 240886 618854
rect 271370 618938 271606 619174
rect 271370 618618 271606 618854
rect 302090 618938 302326 619174
rect 302090 618618 302326 618854
rect 332810 618938 333046 619174
rect 332810 618618 333046 618854
rect 363530 618938 363766 619174
rect 363530 618618 363766 618854
rect 394250 618938 394486 619174
rect 394250 618618 394486 618854
rect 424970 618938 425206 619174
rect 424970 618618 425206 618854
rect 455690 618938 455926 619174
rect 455690 618618 455926 618854
rect 486410 618938 486646 619174
rect 486410 618618 486646 618854
rect 517130 618938 517366 619174
rect 517130 618618 517366 618854
rect 547850 618938 548086 619174
rect 547850 618618 548086 618854
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 10250 615218 10486 615454
rect 10250 614898 10486 615134
rect 40970 615218 41206 615454
rect 40970 614898 41206 615134
rect 71690 615218 71926 615454
rect 71690 614898 71926 615134
rect 102410 615218 102646 615454
rect 102410 614898 102646 615134
rect 133130 615218 133366 615454
rect 133130 614898 133366 615134
rect 163850 615218 164086 615454
rect 163850 614898 164086 615134
rect 194570 615218 194806 615454
rect 194570 614898 194806 615134
rect 225290 615218 225526 615454
rect 225290 614898 225526 615134
rect 256010 615218 256246 615454
rect 256010 614898 256246 615134
rect 286730 615218 286966 615454
rect 286730 614898 286966 615134
rect 317450 615218 317686 615454
rect 317450 614898 317686 615134
rect 348170 615218 348406 615454
rect 348170 614898 348406 615134
rect 378890 615218 379126 615454
rect 378890 614898 379126 615134
rect 409610 615218 409846 615454
rect 409610 614898 409846 615134
rect 440330 615218 440566 615454
rect 440330 614898 440566 615134
rect 471050 615218 471286 615454
rect 471050 614898 471286 615134
rect 501770 615218 502006 615454
rect 501770 614898 502006 615134
rect 532490 615218 532726 615454
rect 532490 614898 532726 615134
rect 563210 615218 563446 615454
rect 563210 614898 563446 615134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 25610 582938 25846 583174
rect 25610 582618 25846 582854
rect 56330 582938 56566 583174
rect 56330 582618 56566 582854
rect 87050 582938 87286 583174
rect 87050 582618 87286 582854
rect 117770 582938 118006 583174
rect 117770 582618 118006 582854
rect 148490 582938 148726 583174
rect 148490 582618 148726 582854
rect 179210 582938 179446 583174
rect 179210 582618 179446 582854
rect 209930 582938 210166 583174
rect 209930 582618 210166 582854
rect 240650 582938 240886 583174
rect 240650 582618 240886 582854
rect 271370 582938 271606 583174
rect 271370 582618 271606 582854
rect 302090 582938 302326 583174
rect 302090 582618 302326 582854
rect 332810 582938 333046 583174
rect 332810 582618 333046 582854
rect 363530 582938 363766 583174
rect 363530 582618 363766 582854
rect 394250 582938 394486 583174
rect 394250 582618 394486 582854
rect 424970 582938 425206 583174
rect 424970 582618 425206 582854
rect 455690 582938 455926 583174
rect 455690 582618 455926 582854
rect 486410 582938 486646 583174
rect 486410 582618 486646 582854
rect 517130 582938 517366 583174
rect 517130 582618 517366 582854
rect 547850 582938 548086 583174
rect 547850 582618 548086 582854
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 10250 579218 10486 579454
rect 10250 578898 10486 579134
rect 40970 579218 41206 579454
rect 40970 578898 41206 579134
rect 71690 579218 71926 579454
rect 71690 578898 71926 579134
rect 102410 579218 102646 579454
rect 102410 578898 102646 579134
rect 133130 579218 133366 579454
rect 133130 578898 133366 579134
rect 163850 579218 164086 579454
rect 163850 578898 164086 579134
rect 194570 579218 194806 579454
rect 194570 578898 194806 579134
rect 225290 579218 225526 579454
rect 225290 578898 225526 579134
rect 256010 579218 256246 579454
rect 256010 578898 256246 579134
rect 286730 579218 286966 579454
rect 286730 578898 286966 579134
rect 317450 579218 317686 579454
rect 317450 578898 317686 579134
rect 348170 579218 348406 579454
rect 348170 578898 348406 579134
rect 378890 579218 379126 579454
rect 378890 578898 379126 579134
rect 409610 579218 409846 579454
rect 409610 578898 409846 579134
rect 440330 579218 440566 579454
rect 440330 578898 440566 579134
rect 471050 579218 471286 579454
rect 471050 578898 471286 579134
rect 501770 579218 502006 579454
rect 501770 578898 502006 579134
rect 532490 579218 532726 579454
rect 532490 578898 532726 579134
rect 563210 579218 563446 579454
rect 563210 578898 563446 579134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 25610 546938 25846 547174
rect 25610 546618 25846 546854
rect 56330 546938 56566 547174
rect 56330 546618 56566 546854
rect 87050 546938 87286 547174
rect 87050 546618 87286 546854
rect 117770 546938 118006 547174
rect 117770 546618 118006 546854
rect 148490 546938 148726 547174
rect 148490 546618 148726 546854
rect 179210 546938 179446 547174
rect 179210 546618 179446 546854
rect 209930 546938 210166 547174
rect 209930 546618 210166 546854
rect 240650 546938 240886 547174
rect 240650 546618 240886 546854
rect 271370 546938 271606 547174
rect 271370 546618 271606 546854
rect 302090 546938 302326 547174
rect 302090 546618 302326 546854
rect 332810 546938 333046 547174
rect 332810 546618 333046 546854
rect 363530 546938 363766 547174
rect 363530 546618 363766 546854
rect 394250 546938 394486 547174
rect 394250 546618 394486 546854
rect 424970 546938 425206 547174
rect 424970 546618 425206 546854
rect 455690 546938 455926 547174
rect 455690 546618 455926 546854
rect 486410 546938 486646 547174
rect 486410 546618 486646 546854
rect 517130 546938 517366 547174
rect 517130 546618 517366 546854
rect 547850 546938 548086 547174
rect 547850 546618 548086 546854
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 10250 543218 10486 543454
rect 10250 542898 10486 543134
rect 40970 543218 41206 543454
rect 40970 542898 41206 543134
rect 71690 543218 71926 543454
rect 71690 542898 71926 543134
rect 102410 543218 102646 543454
rect 102410 542898 102646 543134
rect 133130 543218 133366 543454
rect 133130 542898 133366 543134
rect 163850 543218 164086 543454
rect 163850 542898 164086 543134
rect 194570 543218 194806 543454
rect 194570 542898 194806 543134
rect 225290 543218 225526 543454
rect 225290 542898 225526 543134
rect 256010 543218 256246 543454
rect 256010 542898 256246 543134
rect 286730 543218 286966 543454
rect 286730 542898 286966 543134
rect 317450 543218 317686 543454
rect 317450 542898 317686 543134
rect 348170 543218 348406 543454
rect 348170 542898 348406 543134
rect 378890 543218 379126 543454
rect 378890 542898 379126 543134
rect 409610 543218 409846 543454
rect 409610 542898 409846 543134
rect 440330 543218 440566 543454
rect 440330 542898 440566 543134
rect 471050 543218 471286 543454
rect 471050 542898 471286 543134
rect 501770 543218 502006 543454
rect 501770 542898 502006 543134
rect 532490 543218 532726 543454
rect 532490 542898 532726 543134
rect 563210 543218 563446 543454
rect 563210 542898 563446 543134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 25610 510938 25846 511174
rect 25610 510618 25846 510854
rect 56330 510938 56566 511174
rect 56330 510618 56566 510854
rect 87050 510938 87286 511174
rect 87050 510618 87286 510854
rect 117770 510938 118006 511174
rect 117770 510618 118006 510854
rect 148490 510938 148726 511174
rect 148490 510618 148726 510854
rect 179210 510938 179446 511174
rect 179210 510618 179446 510854
rect 209930 510938 210166 511174
rect 209930 510618 210166 510854
rect 240650 510938 240886 511174
rect 240650 510618 240886 510854
rect 271370 510938 271606 511174
rect 271370 510618 271606 510854
rect 302090 510938 302326 511174
rect 302090 510618 302326 510854
rect 332810 510938 333046 511174
rect 332810 510618 333046 510854
rect 363530 510938 363766 511174
rect 363530 510618 363766 510854
rect 394250 510938 394486 511174
rect 394250 510618 394486 510854
rect 424970 510938 425206 511174
rect 424970 510618 425206 510854
rect 455690 510938 455926 511174
rect 455690 510618 455926 510854
rect 486410 510938 486646 511174
rect 486410 510618 486646 510854
rect 517130 510938 517366 511174
rect 517130 510618 517366 510854
rect 547850 510938 548086 511174
rect 547850 510618 548086 510854
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 10250 507218 10486 507454
rect 10250 506898 10486 507134
rect 40970 507218 41206 507454
rect 40970 506898 41206 507134
rect 71690 507218 71926 507454
rect 71690 506898 71926 507134
rect 102410 507218 102646 507454
rect 102410 506898 102646 507134
rect 133130 507218 133366 507454
rect 133130 506898 133366 507134
rect 163850 507218 164086 507454
rect 163850 506898 164086 507134
rect 194570 507218 194806 507454
rect 194570 506898 194806 507134
rect 225290 507218 225526 507454
rect 225290 506898 225526 507134
rect 256010 507218 256246 507454
rect 256010 506898 256246 507134
rect 286730 507218 286966 507454
rect 286730 506898 286966 507134
rect 317450 507218 317686 507454
rect 317450 506898 317686 507134
rect 348170 507218 348406 507454
rect 348170 506898 348406 507134
rect 378890 507218 379126 507454
rect 378890 506898 379126 507134
rect 409610 507218 409846 507454
rect 409610 506898 409846 507134
rect 440330 507218 440566 507454
rect 440330 506898 440566 507134
rect 471050 507218 471286 507454
rect 471050 506898 471286 507134
rect 501770 507218 502006 507454
rect 501770 506898 502006 507134
rect 532490 507218 532726 507454
rect 532490 506898 532726 507134
rect 563210 507218 563446 507454
rect 563210 506898 563446 507134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 25610 474938 25846 475174
rect 25610 474618 25846 474854
rect 56330 474938 56566 475174
rect 56330 474618 56566 474854
rect 87050 474938 87286 475174
rect 87050 474618 87286 474854
rect 117770 474938 118006 475174
rect 117770 474618 118006 474854
rect 148490 474938 148726 475174
rect 148490 474618 148726 474854
rect 179210 474938 179446 475174
rect 179210 474618 179446 474854
rect 209930 474938 210166 475174
rect 209930 474618 210166 474854
rect 240650 474938 240886 475174
rect 240650 474618 240886 474854
rect 271370 474938 271606 475174
rect 271370 474618 271606 474854
rect 302090 474938 302326 475174
rect 302090 474618 302326 474854
rect 332810 474938 333046 475174
rect 332810 474618 333046 474854
rect 363530 474938 363766 475174
rect 363530 474618 363766 474854
rect 394250 474938 394486 475174
rect 394250 474618 394486 474854
rect 424970 474938 425206 475174
rect 424970 474618 425206 474854
rect 455690 474938 455926 475174
rect 455690 474618 455926 474854
rect 486410 474938 486646 475174
rect 486410 474618 486646 474854
rect 517130 474938 517366 475174
rect 517130 474618 517366 474854
rect 547850 474938 548086 475174
rect 547850 474618 548086 474854
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 10250 471218 10486 471454
rect 10250 470898 10486 471134
rect 40970 471218 41206 471454
rect 40970 470898 41206 471134
rect 71690 471218 71926 471454
rect 71690 470898 71926 471134
rect 102410 471218 102646 471454
rect 102410 470898 102646 471134
rect 133130 471218 133366 471454
rect 133130 470898 133366 471134
rect 163850 471218 164086 471454
rect 163850 470898 164086 471134
rect 194570 471218 194806 471454
rect 194570 470898 194806 471134
rect 225290 471218 225526 471454
rect 225290 470898 225526 471134
rect 256010 471218 256246 471454
rect 256010 470898 256246 471134
rect 286730 471218 286966 471454
rect 286730 470898 286966 471134
rect 317450 471218 317686 471454
rect 317450 470898 317686 471134
rect 348170 471218 348406 471454
rect 348170 470898 348406 471134
rect 378890 471218 379126 471454
rect 378890 470898 379126 471134
rect 409610 471218 409846 471454
rect 409610 470898 409846 471134
rect 440330 471218 440566 471454
rect 440330 470898 440566 471134
rect 471050 471218 471286 471454
rect 471050 470898 471286 471134
rect 501770 471218 502006 471454
rect 501770 470898 502006 471134
rect 532490 471218 532726 471454
rect 532490 470898 532726 471134
rect 563210 471218 563446 471454
rect 563210 470898 563446 471134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 25610 438938 25846 439174
rect 25610 438618 25846 438854
rect 56330 438938 56566 439174
rect 56330 438618 56566 438854
rect 87050 438938 87286 439174
rect 87050 438618 87286 438854
rect 117770 438938 118006 439174
rect 117770 438618 118006 438854
rect 148490 438938 148726 439174
rect 148490 438618 148726 438854
rect 179210 438938 179446 439174
rect 179210 438618 179446 438854
rect 209930 438938 210166 439174
rect 209930 438618 210166 438854
rect 240650 438938 240886 439174
rect 240650 438618 240886 438854
rect 271370 438938 271606 439174
rect 271370 438618 271606 438854
rect 302090 438938 302326 439174
rect 302090 438618 302326 438854
rect 332810 438938 333046 439174
rect 332810 438618 333046 438854
rect 363530 438938 363766 439174
rect 363530 438618 363766 438854
rect 394250 438938 394486 439174
rect 394250 438618 394486 438854
rect 424970 438938 425206 439174
rect 424970 438618 425206 438854
rect 455690 438938 455926 439174
rect 455690 438618 455926 438854
rect 486410 438938 486646 439174
rect 486410 438618 486646 438854
rect 517130 438938 517366 439174
rect 517130 438618 517366 438854
rect 547850 438938 548086 439174
rect 547850 438618 548086 438854
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 10250 435218 10486 435454
rect 10250 434898 10486 435134
rect 40970 435218 41206 435454
rect 40970 434898 41206 435134
rect 71690 435218 71926 435454
rect 71690 434898 71926 435134
rect 102410 435218 102646 435454
rect 102410 434898 102646 435134
rect 133130 435218 133366 435454
rect 133130 434898 133366 435134
rect 163850 435218 164086 435454
rect 163850 434898 164086 435134
rect 194570 435218 194806 435454
rect 194570 434898 194806 435134
rect 225290 435218 225526 435454
rect 225290 434898 225526 435134
rect 256010 435218 256246 435454
rect 256010 434898 256246 435134
rect 286730 435218 286966 435454
rect 286730 434898 286966 435134
rect 317450 435218 317686 435454
rect 317450 434898 317686 435134
rect 348170 435218 348406 435454
rect 348170 434898 348406 435134
rect 378890 435218 379126 435454
rect 378890 434898 379126 435134
rect 409610 435218 409846 435454
rect 409610 434898 409846 435134
rect 440330 435218 440566 435454
rect 440330 434898 440566 435134
rect 471050 435218 471286 435454
rect 471050 434898 471286 435134
rect 501770 435218 502006 435454
rect 501770 434898 502006 435134
rect 532490 435218 532726 435454
rect 532490 434898 532726 435134
rect 563210 435218 563446 435454
rect 563210 434898 563446 435134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 25610 402938 25846 403174
rect 25610 402618 25846 402854
rect 56330 402938 56566 403174
rect 56330 402618 56566 402854
rect 87050 402938 87286 403174
rect 87050 402618 87286 402854
rect 117770 402938 118006 403174
rect 117770 402618 118006 402854
rect 148490 402938 148726 403174
rect 148490 402618 148726 402854
rect 179210 402938 179446 403174
rect 179210 402618 179446 402854
rect 209930 402938 210166 403174
rect 209930 402618 210166 402854
rect 240650 402938 240886 403174
rect 240650 402618 240886 402854
rect 271370 402938 271606 403174
rect 271370 402618 271606 402854
rect 302090 402938 302326 403174
rect 302090 402618 302326 402854
rect 332810 402938 333046 403174
rect 332810 402618 333046 402854
rect 363530 402938 363766 403174
rect 363530 402618 363766 402854
rect 394250 402938 394486 403174
rect 394250 402618 394486 402854
rect 424970 402938 425206 403174
rect 424970 402618 425206 402854
rect 455690 402938 455926 403174
rect 455690 402618 455926 402854
rect 486410 402938 486646 403174
rect 486410 402618 486646 402854
rect 517130 402938 517366 403174
rect 517130 402618 517366 402854
rect 547850 402938 548086 403174
rect 547850 402618 548086 402854
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 10250 399218 10486 399454
rect 10250 398898 10486 399134
rect 40970 399218 41206 399454
rect 40970 398898 41206 399134
rect 71690 399218 71926 399454
rect 71690 398898 71926 399134
rect 102410 399218 102646 399454
rect 102410 398898 102646 399134
rect 133130 399218 133366 399454
rect 133130 398898 133366 399134
rect 163850 399218 164086 399454
rect 163850 398898 164086 399134
rect 194570 399218 194806 399454
rect 194570 398898 194806 399134
rect 225290 399218 225526 399454
rect 225290 398898 225526 399134
rect 256010 399218 256246 399454
rect 256010 398898 256246 399134
rect 286730 399218 286966 399454
rect 286730 398898 286966 399134
rect 317450 399218 317686 399454
rect 317450 398898 317686 399134
rect 348170 399218 348406 399454
rect 348170 398898 348406 399134
rect 378890 399218 379126 399454
rect 378890 398898 379126 399134
rect 409610 399218 409846 399454
rect 409610 398898 409846 399134
rect 440330 399218 440566 399454
rect 440330 398898 440566 399134
rect 471050 399218 471286 399454
rect 471050 398898 471286 399134
rect 501770 399218 502006 399454
rect 501770 398898 502006 399134
rect 532490 399218 532726 399454
rect 532490 398898 532726 399134
rect 563210 399218 563446 399454
rect 563210 398898 563446 399134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 25610 366938 25846 367174
rect 25610 366618 25846 366854
rect 56330 366938 56566 367174
rect 56330 366618 56566 366854
rect 87050 366938 87286 367174
rect 87050 366618 87286 366854
rect 117770 366938 118006 367174
rect 117770 366618 118006 366854
rect 148490 366938 148726 367174
rect 148490 366618 148726 366854
rect 179210 366938 179446 367174
rect 179210 366618 179446 366854
rect 209930 366938 210166 367174
rect 209930 366618 210166 366854
rect 240650 366938 240886 367174
rect 240650 366618 240886 366854
rect 271370 366938 271606 367174
rect 271370 366618 271606 366854
rect 302090 366938 302326 367174
rect 302090 366618 302326 366854
rect 332810 366938 333046 367174
rect 332810 366618 333046 366854
rect 363530 366938 363766 367174
rect 363530 366618 363766 366854
rect 394250 366938 394486 367174
rect 394250 366618 394486 366854
rect 424970 366938 425206 367174
rect 424970 366618 425206 366854
rect 455690 366938 455926 367174
rect 455690 366618 455926 366854
rect 486410 366938 486646 367174
rect 486410 366618 486646 366854
rect 517130 366938 517366 367174
rect 517130 366618 517366 366854
rect 547850 366938 548086 367174
rect 547850 366618 548086 366854
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 10250 363218 10486 363454
rect 10250 362898 10486 363134
rect 40970 363218 41206 363454
rect 40970 362898 41206 363134
rect 71690 363218 71926 363454
rect 71690 362898 71926 363134
rect 102410 363218 102646 363454
rect 102410 362898 102646 363134
rect 133130 363218 133366 363454
rect 133130 362898 133366 363134
rect 163850 363218 164086 363454
rect 163850 362898 164086 363134
rect 194570 363218 194806 363454
rect 194570 362898 194806 363134
rect 225290 363218 225526 363454
rect 225290 362898 225526 363134
rect 256010 363218 256246 363454
rect 256010 362898 256246 363134
rect 286730 363218 286966 363454
rect 286730 362898 286966 363134
rect 317450 363218 317686 363454
rect 317450 362898 317686 363134
rect 348170 363218 348406 363454
rect 348170 362898 348406 363134
rect 378890 363218 379126 363454
rect 378890 362898 379126 363134
rect 409610 363218 409846 363454
rect 409610 362898 409846 363134
rect 440330 363218 440566 363454
rect 440330 362898 440566 363134
rect 471050 363218 471286 363454
rect 471050 362898 471286 363134
rect 501770 363218 502006 363454
rect 501770 362898 502006 363134
rect 532490 363218 532726 363454
rect 532490 362898 532726 363134
rect 563210 363218 563446 363454
rect 563210 362898 563446 363134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 25610 330938 25846 331174
rect 25610 330618 25846 330854
rect 56330 330938 56566 331174
rect 56330 330618 56566 330854
rect 87050 330938 87286 331174
rect 87050 330618 87286 330854
rect 117770 330938 118006 331174
rect 117770 330618 118006 330854
rect 148490 330938 148726 331174
rect 148490 330618 148726 330854
rect 179210 330938 179446 331174
rect 179210 330618 179446 330854
rect 209930 330938 210166 331174
rect 209930 330618 210166 330854
rect 240650 330938 240886 331174
rect 240650 330618 240886 330854
rect 271370 330938 271606 331174
rect 271370 330618 271606 330854
rect 302090 330938 302326 331174
rect 302090 330618 302326 330854
rect 332810 330938 333046 331174
rect 332810 330618 333046 330854
rect 363530 330938 363766 331174
rect 363530 330618 363766 330854
rect 394250 330938 394486 331174
rect 394250 330618 394486 330854
rect 424970 330938 425206 331174
rect 424970 330618 425206 330854
rect 455690 330938 455926 331174
rect 455690 330618 455926 330854
rect 486410 330938 486646 331174
rect 486410 330618 486646 330854
rect 517130 330938 517366 331174
rect 517130 330618 517366 330854
rect 547850 330938 548086 331174
rect 547850 330618 548086 330854
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 10250 327218 10486 327454
rect 10250 326898 10486 327134
rect 40970 327218 41206 327454
rect 40970 326898 41206 327134
rect 71690 327218 71926 327454
rect 71690 326898 71926 327134
rect 102410 327218 102646 327454
rect 102410 326898 102646 327134
rect 133130 327218 133366 327454
rect 133130 326898 133366 327134
rect 163850 327218 164086 327454
rect 163850 326898 164086 327134
rect 194570 327218 194806 327454
rect 194570 326898 194806 327134
rect 225290 327218 225526 327454
rect 225290 326898 225526 327134
rect 256010 327218 256246 327454
rect 256010 326898 256246 327134
rect 286730 327218 286966 327454
rect 286730 326898 286966 327134
rect 317450 327218 317686 327454
rect 317450 326898 317686 327134
rect 348170 327218 348406 327454
rect 348170 326898 348406 327134
rect 378890 327218 379126 327454
rect 378890 326898 379126 327134
rect 409610 327218 409846 327454
rect 409610 326898 409846 327134
rect 440330 327218 440566 327454
rect 440330 326898 440566 327134
rect 471050 327218 471286 327454
rect 471050 326898 471286 327134
rect 501770 327218 502006 327454
rect 501770 326898 502006 327134
rect 532490 327218 532726 327454
rect 532490 326898 532726 327134
rect 563210 327218 563446 327454
rect 563210 326898 563446 327134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 25610 294938 25846 295174
rect 25610 294618 25846 294854
rect 56330 294938 56566 295174
rect 56330 294618 56566 294854
rect 87050 294938 87286 295174
rect 87050 294618 87286 294854
rect 117770 294938 118006 295174
rect 117770 294618 118006 294854
rect 148490 294938 148726 295174
rect 148490 294618 148726 294854
rect 179210 294938 179446 295174
rect 179210 294618 179446 294854
rect 209930 294938 210166 295174
rect 209930 294618 210166 294854
rect 240650 294938 240886 295174
rect 240650 294618 240886 294854
rect 271370 294938 271606 295174
rect 271370 294618 271606 294854
rect 302090 294938 302326 295174
rect 302090 294618 302326 294854
rect 332810 294938 333046 295174
rect 332810 294618 333046 294854
rect 363530 294938 363766 295174
rect 363530 294618 363766 294854
rect 394250 294938 394486 295174
rect 394250 294618 394486 294854
rect 424970 294938 425206 295174
rect 424970 294618 425206 294854
rect 455690 294938 455926 295174
rect 455690 294618 455926 294854
rect 486410 294938 486646 295174
rect 486410 294618 486646 294854
rect 517130 294938 517366 295174
rect 517130 294618 517366 294854
rect 547850 294938 548086 295174
rect 547850 294618 548086 294854
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 10250 291218 10486 291454
rect 10250 290898 10486 291134
rect 40970 291218 41206 291454
rect 40970 290898 41206 291134
rect 71690 291218 71926 291454
rect 71690 290898 71926 291134
rect 102410 291218 102646 291454
rect 102410 290898 102646 291134
rect 133130 291218 133366 291454
rect 133130 290898 133366 291134
rect 163850 291218 164086 291454
rect 163850 290898 164086 291134
rect 194570 291218 194806 291454
rect 194570 290898 194806 291134
rect 225290 291218 225526 291454
rect 225290 290898 225526 291134
rect 256010 291218 256246 291454
rect 256010 290898 256246 291134
rect 286730 291218 286966 291454
rect 286730 290898 286966 291134
rect 317450 291218 317686 291454
rect 317450 290898 317686 291134
rect 348170 291218 348406 291454
rect 348170 290898 348406 291134
rect 378890 291218 379126 291454
rect 378890 290898 379126 291134
rect 409610 291218 409846 291454
rect 409610 290898 409846 291134
rect 440330 291218 440566 291454
rect 440330 290898 440566 291134
rect 471050 291218 471286 291454
rect 471050 290898 471286 291134
rect 501770 291218 502006 291454
rect 501770 290898 502006 291134
rect 532490 291218 532726 291454
rect 532490 290898 532726 291134
rect 563210 291218 563446 291454
rect 563210 290898 563446 291134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 25610 258938 25846 259174
rect 25610 258618 25846 258854
rect 56330 258938 56566 259174
rect 56330 258618 56566 258854
rect 87050 258938 87286 259174
rect 87050 258618 87286 258854
rect 117770 258938 118006 259174
rect 117770 258618 118006 258854
rect 148490 258938 148726 259174
rect 148490 258618 148726 258854
rect 179210 258938 179446 259174
rect 179210 258618 179446 258854
rect 209930 258938 210166 259174
rect 209930 258618 210166 258854
rect 240650 258938 240886 259174
rect 240650 258618 240886 258854
rect 271370 258938 271606 259174
rect 271370 258618 271606 258854
rect 302090 258938 302326 259174
rect 302090 258618 302326 258854
rect 332810 258938 333046 259174
rect 332810 258618 333046 258854
rect 363530 258938 363766 259174
rect 363530 258618 363766 258854
rect 394250 258938 394486 259174
rect 394250 258618 394486 258854
rect 424970 258938 425206 259174
rect 424970 258618 425206 258854
rect 455690 258938 455926 259174
rect 455690 258618 455926 258854
rect 486410 258938 486646 259174
rect 486410 258618 486646 258854
rect 517130 258938 517366 259174
rect 517130 258618 517366 258854
rect 547850 258938 548086 259174
rect 547850 258618 548086 258854
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 10250 255218 10486 255454
rect 10250 254898 10486 255134
rect 40970 255218 41206 255454
rect 40970 254898 41206 255134
rect 71690 255218 71926 255454
rect 71690 254898 71926 255134
rect 102410 255218 102646 255454
rect 102410 254898 102646 255134
rect 133130 255218 133366 255454
rect 133130 254898 133366 255134
rect 163850 255218 164086 255454
rect 163850 254898 164086 255134
rect 194570 255218 194806 255454
rect 194570 254898 194806 255134
rect 225290 255218 225526 255454
rect 225290 254898 225526 255134
rect 256010 255218 256246 255454
rect 256010 254898 256246 255134
rect 286730 255218 286966 255454
rect 286730 254898 286966 255134
rect 317450 255218 317686 255454
rect 317450 254898 317686 255134
rect 348170 255218 348406 255454
rect 348170 254898 348406 255134
rect 378890 255218 379126 255454
rect 378890 254898 379126 255134
rect 409610 255218 409846 255454
rect 409610 254898 409846 255134
rect 440330 255218 440566 255454
rect 440330 254898 440566 255134
rect 471050 255218 471286 255454
rect 471050 254898 471286 255134
rect 501770 255218 502006 255454
rect 501770 254898 502006 255134
rect 532490 255218 532726 255454
rect 532490 254898 532726 255134
rect 563210 255218 563446 255454
rect 563210 254898 563446 255134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 25610 222938 25846 223174
rect 25610 222618 25846 222854
rect 56330 222938 56566 223174
rect 56330 222618 56566 222854
rect 87050 222938 87286 223174
rect 87050 222618 87286 222854
rect 117770 222938 118006 223174
rect 117770 222618 118006 222854
rect 148490 222938 148726 223174
rect 148490 222618 148726 222854
rect 179210 222938 179446 223174
rect 179210 222618 179446 222854
rect 209930 222938 210166 223174
rect 209930 222618 210166 222854
rect 240650 222938 240886 223174
rect 240650 222618 240886 222854
rect 271370 222938 271606 223174
rect 271370 222618 271606 222854
rect 302090 222938 302326 223174
rect 302090 222618 302326 222854
rect 332810 222938 333046 223174
rect 332810 222618 333046 222854
rect 363530 222938 363766 223174
rect 363530 222618 363766 222854
rect 394250 222938 394486 223174
rect 394250 222618 394486 222854
rect 424970 222938 425206 223174
rect 424970 222618 425206 222854
rect 455690 222938 455926 223174
rect 455690 222618 455926 222854
rect 486410 222938 486646 223174
rect 486410 222618 486646 222854
rect 517130 222938 517366 223174
rect 517130 222618 517366 222854
rect 547850 222938 548086 223174
rect 547850 222618 548086 222854
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 10250 219218 10486 219454
rect 10250 218898 10486 219134
rect 40970 219218 41206 219454
rect 40970 218898 41206 219134
rect 71690 219218 71926 219454
rect 71690 218898 71926 219134
rect 102410 219218 102646 219454
rect 102410 218898 102646 219134
rect 133130 219218 133366 219454
rect 133130 218898 133366 219134
rect 163850 219218 164086 219454
rect 163850 218898 164086 219134
rect 194570 219218 194806 219454
rect 194570 218898 194806 219134
rect 225290 219218 225526 219454
rect 225290 218898 225526 219134
rect 256010 219218 256246 219454
rect 256010 218898 256246 219134
rect 286730 219218 286966 219454
rect 286730 218898 286966 219134
rect 317450 219218 317686 219454
rect 317450 218898 317686 219134
rect 348170 219218 348406 219454
rect 348170 218898 348406 219134
rect 378890 219218 379126 219454
rect 378890 218898 379126 219134
rect 409610 219218 409846 219454
rect 409610 218898 409846 219134
rect 440330 219218 440566 219454
rect 440330 218898 440566 219134
rect 471050 219218 471286 219454
rect 471050 218898 471286 219134
rect 501770 219218 502006 219454
rect 501770 218898 502006 219134
rect 532490 219218 532726 219454
rect 532490 218898 532726 219134
rect 563210 219218 563446 219454
rect 563210 218898 563446 219134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 25610 186938 25846 187174
rect 25610 186618 25846 186854
rect 56330 186938 56566 187174
rect 56330 186618 56566 186854
rect 87050 186938 87286 187174
rect 87050 186618 87286 186854
rect 117770 186938 118006 187174
rect 117770 186618 118006 186854
rect 148490 186938 148726 187174
rect 148490 186618 148726 186854
rect 179210 186938 179446 187174
rect 179210 186618 179446 186854
rect 209930 186938 210166 187174
rect 209930 186618 210166 186854
rect 240650 186938 240886 187174
rect 240650 186618 240886 186854
rect 271370 186938 271606 187174
rect 271370 186618 271606 186854
rect 302090 186938 302326 187174
rect 302090 186618 302326 186854
rect 332810 186938 333046 187174
rect 332810 186618 333046 186854
rect 363530 186938 363766 187174
rect 363530 186618 363766 186854
rect 394250 186938 394486 187174
rect 394250 186618 394486 186854
rect 424970 186938 425206 187174
rect 424970 186618 425206 186854
rect 455690 186938 455926 187174
rect 455690 186618 455926 186854
rect 486410 186938 486646 187174
rect 486410 186618 486646 186854
rect 517130 186938 517366 187174
rect 517130 186618 517366 186854
rect 547850 186938 548086 187174
rect 547850 186618 548086 186854
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 10250 183218 10486 183454
rect 10250 182898 10486 183134
rect 40970 183218 41206 183454
rect 40970 182898 41206 183134
rect 71690 183218 71926 183454
rect 71690 182898 71926 183134
rect 102410 183218 102646 183454
rect 102410 182898 102646 183134
rect 133130 183218 133366 183454
rect 133130 182898 133366 183134
rect 163850 183218 164086 183454
rect 163850 182898 164086 183134
rect 194570 183218 194806 183454
rect 194570 182898 194806 183134
rect 225290 183218 225526 183454
rect 225290 182898 225526 183134
rect 256010 183218 256246 183454
rect 256010 182898 256246 183134
rect 286730 183218 286966 183454
rect 286730 182898 286966 183134
rect 317450 183218 317686 183454
rect 317450 182898 317686 183134
rect 348170 183218 348406 183454
rect 348170 182898 348406 183134
rect 378890 183218 379126 183454
rect 378890 182898 379126 183134
rect 409610 183218 409846 183454
rect 409610 182898 409846 183134
rect 440330 183218 440566 183454
rect 440330 182898 440566 183134
rect 471050 183218 471286 183454
rect 471050 182898 471286 183134
rect 501770 183218 502006 183454
rect 501770 182898 502006 183134
rect 532490 183218 532726 183454
rect 532490 182898 532726 183134
rect 563210 183218 563446 183454
rect 563210 182898 563446 183134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 25610 150938 25846 151174
rect 25610 150618 25846 150854
rect 56330 150938 56566 151174
rect 56330 150618 56566 150854
rect 87050 150938 87286 151174
rect 87050 150618 87286 150854
rect 117770 150938 118006 151174
rect 117770 150618 118006 150854
rect 148490 150938 148726 151174
rect 148490 150618 148726 150854
rect 179210 150938 179446 151174
rect 179210 150618 179446 150854
rect 209930 150938 210166 151174
rect 209930 150618 210166 150854
rect 240650 150938 240886 151174
rect 240650 150618 240886 150854
rect 271370 150938 271606 151174
rect 271370 150618 271606 150854
rect 302090 150938 302326 151174
rect 302090 150618 302326 150854
rect 332810 150938 333046 151174
rect 332810 150618 333046 150854
rect 363530 150938 363766 151174
rect 363530 150618 363766 150854
rect 394250 150938 394486 151174
rect 394250 150618 394486 150854
rect 424970 150938 425206 151174
rect 424970 150618 425206 150854
rect 455690 150938 455926 151174
rect 455690 150618 455926 150854
rect 486410 150938 486646 151174
rect 486410 150618 486646 150854
rect 517130 150938 517366 151174
rect 517130 150618 517366 150854
rect 547850 150938 548086 151174
rect 547850 150618 548086 150854
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 10250 147218 10486 147454
rect 10250 146898 10486 147134
rect 40970 147218 41206 147454
rect 40970 146898 41206 147134
rect 71690 147218 71926 147454
rect 71690 146898 71926 147134
rect 102410 147218 102646 147454
rect 102410 146898 102646 147134
rect 133130 147218 133366 147454
rect 133130 146898 133366 147134
rect 163850 147218 164086 147454
rect 163850 146898 164086 147134
rect 194570 147218 194806 147454
rect 194570 146898 194806 147134
rect 225290 147218 225526 147454
rect 225290 146898 225526 147134
rect 256010 147218 256246 147454
rect 256010 146898 256246 147134
rect 286730 147218 286966 147454
rect 286730 146898 286966 147134
rect 317450 147218 317686 147454
rect 317450 146898 317686 147134
rect 348170 147218 348406 147454
rect 348170 146898 348406 147134
rect 378890 147218 379126 147454
rect 378890 146898 379126 147134
rect 409610 147218 409846 147454
rect 409610 146898 409846 147134
rect 440330 147218 440566 147454
rect 440330 146898 440566 147134
rect 471050 147218 471286 147454
rect 471050 146898 471286 147134
rect 501770 147218 502006 147454
rect 501770 146898 502006 147134
rect 532490 147218 532726 147454
rect 532490 146898 532726 147134
rect 563210 147218 563446 147454
rect 563210 146898 563446 147134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 25610 114938 25846 115174
rect 25610 114618 25846 114854
rect 56330 114938 56566 115174
rect 56330 114618 56566 114854
rect 87050 114938 87286 115174
rect 87050 114618 87286 114854
rect 117770 114938 118006 115174
rect 117770 114618 118006 114854
rect 148490 114938 148726 115174
rect 148490 114618 148726 114854
rect 179210 114938 179446 115174
rect 179210 114618 179446 114854
rect 209930 114938 210166 115174
rect 209930 114618 210166 114854
rect 240650 114938 240886 115174
rect 240650 114618 240886 114854
rect 271370 114938 271606 115174
rect 271370 114618 271606 114854
rect 302090 114938 302326 115174
rect 302090 114618 302326 114854
rect 332810 114938 333046 115174
rect 332810 114618 333046 114854
rect 363530 114938 363766 115174
rect 363530 114618 363766 114854
rect 394250 114938 394486 115174
rect 394250 114618 394486 114854
rect 424970 114938 425206 115174
rect 424970 114618 425206 114854
rect 455690 114938 455926 115174
rect 455690 114618 455926 114854
rect 486410 114938 486646 115174
rect 486410 114618 486646 114854
rect 517130 114938 517366 115174
rect 517130 114618 517366 114854
rect 547850 114938 548086 115174
rect 547850 114618 548086 114854
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 10250 111218 10486 111454
rect 10250 110898 10486 111134
rect 40970 111218 41206 111454
rect 40970 110898 41206 111134
rect 71690 111218 71926 111454
rect 71690 110898 71926 111134
rect 102410 111218 102646 111454
rect 102410 110898 102646 111134
rect 133130 111218 133366 111454
rect 133130 110898 133366 111134
rect 163850 111218 164086 111454
rect 163850 110898 164086 111134
rect 194570 111218 194806 111454
rect 194570 110898 194806 111134
rect 225290 111218 225526 111454
rect 225290 110898 225526 111134
rect 256010 111218 256246 111454
rect 256010 110898 256246 111134
rect 286730 111218 286966 111454
rect 286730 110898 286966 111134
rect 317450 111218 317686 111454
rect 317450 110898 317686 111134
rect 348170 111218 348406 111454
rect 348170 110898 348406 111134
rect 378890 111218 379126 111454
rect 378890 110898 379126 111134
rect 409610 111218 409846 111454
rect 409610 110898 409846 111134
rect 440330 111218 440566 111454
rect 440330 110898 440566 111134
rect 471050 111218 471286 111454
rect 471050 110898 471286 111134
rect 501770 111218 502006 111454
rect 501770 110898 502006 111134
rect 532490 111218 532726 111454
rect 532490 110898 532726 111134
rect 563210 111218 563446 111454
rect 563210 110898 563446 111134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 25610 78938 25846 79174
rect 25610 78618 25846 78854
rect 56330 78938 56566 79174
rect 56330 78618 56566 78854
rect 87050 78938 87286 79174
rect 87050 78618 87286 78854
rect 117770 78938 118006 79174
rect 117770 78618 118006 78854
rect 148490 78938 148726 79174
rect 148490 78618 148726 78854
rect 179210 78938 179446 79174
rect 179210 78618 179446 78854
rect 209930 78938 210166 79174
rect 209930 78618 210166 78854
rect 240650 78938 240886 79174
rect 240650 78618 240886 78854
rect 271370 78938 271606 79174
rect 271370 78618 271606 78854
rect 302090 78938 302326 79174
rect 302090 78618 302326 78854
rect 332810 78938 333046 79174
rect 332810 78618 333046 78854
rect 363530 78938 363766 79174
rect 363530 78618 363766 78854
rect 394250 78938 394486 79174
rect 394250 78618 394486 78854
rect 424970 78938 425206 79174
rect 424970 78618 425206 78854
rect 455690 78938 455926 79174
rect 455690 78618 455926 78854
rect 486410 78938 486646 79174
rect 486410 78618 486646 78854
rect 517130 78938 517366 79174
rect 517130 78618 517366 78854
rect 547850 78938 548086 79174
rect 547850 78618 548086 78854
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 10250 75218 10486 75454
rect 10250 74898 10486 75134
rect 40970 75218 41206 75454
rect 40970 74898 41206 75134
rect 71690 75218 71926 75454
rect 71690 74898 71926 75134
rect 102410 75218 102646 75454
rect 102410 74898 102646 75134
rect 133130 75218 133366 75454
rect 133130 74898 133366 75134
rect 163850 75218 164086 75454
rect 163850 74898 164086 75134
rect 194570 75218 194806 75454
rect 194570 74898 194806 75134
rect 225290 75218 225526 75454
rect 225290 74898 225526 75134
rect 256010 75218 256246 75454
rect 256010 74898 256246 75134
rect 286730 75218 286966 75454
rect 286730 74898 286966 75134
rect 317450 75218 317686 75454
rect 317450 74898 317686 75134
rect 348170 75218 348406 75454
rect 348170 74898 348406 75134
rect 378890 75218 379126 75454
rect 378890 74898 379126 75134
rect 409610 75218 409846 75454
rect 409610 74898 409846 75134
rect 440330 75218 440566 75454
rect 440330 74898 440566 75134
rect 471050 75218 471286 75454
rect 471050 74898 471286 75134
rect 501770 75218 502006 75454
rect 501770 74898 502006 75134
rect 532490 75218 532726 75454
rect 532490 74898 532726 75134
rect 563210 75218 563446 75454
rect 563210 74898 563446 75134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 25610 42938 25846 43174
rect 25610 42618 25846 42854
rect 56330 42938 56566 43174
rect 56330 42618 56566 42854
rect 87050 42938 87286 43174
rect 87050 42618 87286 42854
rect 117770 42938 118006 43174
rect 117770 42618 118006 42854
rect 148490 42938 148726 43174
rect 148490 42618 148726 42854
rect 179210 42938 179446 43174
rect 179210 42618 179446 42854
rect 209930 42938 210166 43174
rect 209930 42618 210166 42854
rect 240650 42938 240886 43174
rect 240650 42618 240886 42854
rect 271370 42938 271606 43174
rect 271370 42618 271606 42854
rect 302090 42938 302326 43174
rect 302090 42618 302326 42854
rect 332810 42938 333046 43174
rect 332810 42618 333046 42854
rect 363530 42938 363766 43174
rect 363530 42618 363766 42854
rect 394250 42938 394486 43174
rect 394250 42618 394486 42854
rect 424970 42938 425206 43174
rect 424970 42618 425206 42854
rect 455690 42938 455926 43174
rect 455690 42618 455926 42854
rect 486410 42938 486646 43174
rect 486410 42618 486646 42854
rect 517130 42938 517366 43174
rect 517130 42618 517366 42854
rect 547850 42938 548086 43174
rect 547850 42618 548086 42854
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 10250 39218 10486 39454
rect 10250 38898 10486 39134
rect 40970 39218 41206 39454
rect 40970 38898 41206 39134
rect 71690 39218 71926 39454
rect 71690 38898 71926 39134
rect 102410 39218 102646 39454
rect 102410 38898 102646 39134
rect 133130 39218 133366 39454
rect 133130 38898 133366 39134
rect 163850 39218 164086 39454
rect 163850 38898 164086 39134
rect 194570 39218 194806 39454
rect 194570 38898 194806 39134
rect 225290 39218 225526 39454
rect 225290 38898 225526 39134
rect 256010 39218 256246 39454
rect 256010 38898 256246 39134
rect 286730 39218 286966 39454
rect 286730 38898 286966 39134
rect 317450 39218 317686 39454
rect 317450 38898 317686 39134
rect 348170 39218 348406 39454
rect 348170 38898 348406 39134
rect 378890 39218 379126 39454
rect 378890 38898 379126 39134
rect 409610 39218 409846 39454
rect 409610 38898 409846 39134
rect 440330 39218 440566 39454
rect 440330 38898 440566 39134
rect 471050 39218 471286 39454
rect 471050 38898 471286 39134
rect 501770 39218 502006 39454
rect 501770 38898 502006 39134
rect 532490 39218 532726 39454
rect 532490 38898 532726 39134
rect 563210 39218 563446 39454
rect 563210 38898 563446 39134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect 5546 -1542 5782 -1306
rect 5866 -1542 6102 -1306
rect 5546 -1862 5782 -1626
rect 5866 -1862 6102 -1626
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -1542 41782 -1306
rect 41866 -1542 42102 -1306
rect 41546 -1862 41782 -1626
rect 41866 -1862 42102 -1626
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -1542 77782 -1306
rect 77866 -1542 78102 -1306
rect 77546 -1862 77782 -1626
rect 77866 -1862 78102 -1626
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -1542 113782 -1306
rect 113866 -1542 114102 -1306
rect 113546 -1862 113782 -1626
rect 113866 -1862 114102 -1626
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -1542 149782 -1306
rect 149866 -1542 150102 -1306
rect 149546 -1862 149782 -1626
rect 149866 -1862 150102 -1626
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -1542 185782 -1306
rect 185866 -1542 186102 -1306
rect 185546 -1862 185782 -1626
rect 185866 -1862 186102 -1626
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -1542 221782 -1306
rect 221866 -1542 222102 -1306
rect 221546 -1862 221782 -1626
rect 221866 -1862 222102 -1626
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -1542 257782 -1306
rect 257866 -1542 258102 -1306
rect 257546 -1862 257782 -1626
rect 257866 -1862 258102 -1626
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -1542 293782 -1306
rect 293866 -1542 294102 -1306
rect 293546 -1862 293782 -1626
rect 293866 -1862 294102 -1626
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -1542 329782 -1306
rect 329866 -1542 330102 -1306
rect 329546 -1862 329782 -1626
rect 329866 -1862 330102 -1626
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -1542 365782 -1306
rect 365866 -1542 366102 -1306
rect 365546 -1862 365782 -1626
rect 365866 -1862 366102 -1626
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -1542 401782 -1306
rect 401866 -1542 402102 -1306
rect 401546 -1862 401782 -1626
rect 401866 -1862 402102 -1626
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -1542 437782 -1306
rect 437866 -1542 438102 -1306
rect 437546 -1862 437782 -1626
rect 437866 -1862 438102 -1626
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -1542 473782 -1306
rect 473866 -1542 474102 -1306
rect 473546 -1862 473782 -1626
rect 473866 -1862 474102 -1626
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -1542 509782 -1306
rect 509866 -1542 510102 -1306
rect 509546 -1862 509782 -1626
rect 509866 -1862 510102 -1626
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -1542 545782 -1306
rect 545866 -1542 546102 -1306
rect 545546 -1862 545782 -1626
rect 545866 -1862 546102 -1626
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 581546 705562 581782 705798
rect 581866 705562 582102 705798
rect 581546 705242 581782 705478
rect 581866 705242 582102 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 690938 586538 691174
rect 586622 690938 586858 691174
rect 586302 690618 586538 690854
rect 586622 690618 586858 690854
rect 586302 654938 586538 655174
rect 586622 654938 586858 655174
rect 586302 654618 586538 654854
rect 586622 654618 586858 654854
rect 586302 618938 586538 619174
rect 586622 618938 586858 619174
rect 586302 618618 586538 618854
rect 586622 618618 586858 618854
rect 586302 582938 586538 583174
rect 586622 582938 586858 583174
rect 586302 582618 586538 582854
rect 586622 582618 586858 582854
rect 586302 546938 586538 547174
rect 586622 546938 586858 547174
rect 586302 546618 586538 546854
rect 586622 546618 586858 546854
rect 586302 510938 586538 511174
rect 586622 510938 586858 511174
rect 586302 510618 586538 510854
rect 586622 510618 586858 510854
rect 586302 474938 586538 475174
rect 586622 474938 586858 475174
rect 586302 474618 586538 474854
rect 586622 474618 586858 474854
rect 586302 438938 586538 439174
rect 586622 438938 586858 439174
rect 586302 438618 586538 438854
rect 586622 438618 586858 438854
rect 586302 402938 586538 403174
rect 586622 402938 586858 403174
rect 586302 402618 586538 402854
rect 586622 402618 586858 402854
rect 586302 366938 586538 367174
rect 586622 366938 586858 367174
rect 586302 366618 586538 366854
rect 586622 366618 586858 366854
rect 586302 330938 586538 331174
rect 586622 330938 586858 331174
rect 586302 330618 586538 330854
rect 586622 330618 586858 330854
rect 586302 294938 586538 295174
rect 586622 294938 586858 295174
rect 586302 294618 586538 294854
rect 586622 294618 586858 294854
rect 586302 258938 586538 259174
rect 586622 258938 586858 259174
rect 586302 258618 586538 258854
rect 586622 258618 586858 258854
rect 586302 222938 586538 223174
rect 586622 222938 586858 223174
rect 586302 222618 586538 222854
rect 586622 222618 586858 222854
rect 586302 186938 586538 187174
rect 586622 186938 586858 187174
rect 586302 186618 586538 186854
rect 586622 186618 586858 186854
rect 586302 150938 586538 151174
rect 586622 150938 586858 151174
rect 586302 150618 586538 150854
rect 586622 150618 586858 150854
rect 586302 114938 586538 115174
rect 586622 114938 586858 115174
rect 586302 114618 586538 114854
rect 586622 114618 586858 114854
rect 586302 78938 586538 79174
rect 586622 78938 586858 79174
rect 586302 78618 586538 78854
rect 586622 78618 586858 78854
rect 586302 42938 586538 43174
rect 586622 42938 586858 43174
rect 586302 42618 586538 42854
rect 586622 42618 586858 42854
rect 586302 6938 586538 7174
rect 586622 6938 586858 7174
rect 586302 6618 586538 6854
rect 586622 6618 586858 6854
rect 581546 -1542 581782 -1306
rect 581866 -1542 582102 -1306
rect 581546 -1862 581782 -1626
rect 581866 -1862 582102 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 694658 587498 694894
rect 587582 694658 587818 694894
rect 587262 694338 587498 694574
rect 587582 694338 587818 694574
rect 587262 658658 587498 658894
rect 587582 658658 587818 658894
rect 587262 658338 587498 658574
rect 587582 658338 587818 658574
rect 587262 622658 587498 622894
rect 587582 622658 587818 622894
rect 587262 622338 587498 622574
rect 587582 622338 587818 622574
rect 587262 586658 587498 586894
rect 587582 586658 587818 586894
rect 587262 586338 587498 586574
rect 587582 586338 587818 586574
rect 587262 550658 587498 550894
rect 587582 550658 587818 550894
rect 587262 550338 587498 550574
rect 587582 550338 587818 550574
rect 587262 514658 587498 514894
rect 587582 514658 587818 514894
rect 587262 514338 587498 514574
rect 587582 514338 587818 514574
rect 587262 478658 587498 478894
rect 587582 478658 587818 478894
rect 587262 478338 587498 478574
rect 587582 478338 587818 478574
rect 587262 442658 587498 442894
rect 587582 442658 587818 442894
rect 587262 442338 587498 442574
rect 587582 442338 587818 442574
rect 587262 406658 587498 406894
rect 587582 406658 587818 406894
rect 587262 406338 587498 406574
rect 587582 406338 587818 406574
rect 587262 370658 587498 370894
rect 587582 370658 587818 370894
rect 587262 370338 587498 370574
rect 587582 370338 587818 370574
rect 587262 334658 587498 334894
rect 587582 334658 587818 334894
rect 587262 334338 587498 334574
rect 587582 334338 587818 334574
rect 587262 298658 587498 298894
rect 587582 298658 587818 298894
rect 587262 298338 587498 298574
rect 587582 298338 587818 298574
rect 587262 262658 587498 262894
rect 587582 262658 587818 262894
rect 587262 262338 587498 262574
rect 587582 262338 587818 262574
rect 587262 226658 587498 226894
rect 587582 226658 587818 226894
rect 587262 226338 587498 226574
rect 587582 226338 587818 226574
rect 587262 190658 587498 190894
rect 587582 190658 587818 190894
rect 587262 190338 587498 190574
rect 587582 190338 587818 190574
rect 587262 154658 587498 154894
rect 587582 154658 587818 154894
rect 587262 154338 587498 154574
rect 587582 154338 587818 154574
rect 587262 118658 587498 118894
rect 587582 118658 587818 118894
rect 587262 118338 587498 118574
rect 587582 118338 587818 118574
rect 587262 82658 587498 82894
rect 587582 82658 587818 82894
rect 587262 82338 587498 82574
rect 587582 82338 587818 82574
rect 587262 46658 587498 46894
rect 587582 46658 587818 46894
rect 587262 46338 587498 46574
rect 587582 46338 587818 46574
rect 587262 10658 587498 10894
rect 587582 10658 587818 10894
rect 587262 10338 587498 10574
rect 587582 10338 587818 10574
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 698378 588458 698614
rect 588542 698378 588778 698614
rect 588222 698058 588458 698294
rect 588542 698058 588778 698294
rect 588222 662378 588458 662614
rect 588542 662378 588778 662614
rect 588222 662058 588458 662294
rect 588542 662058 588778 662294
rect 588222 626378 588458 626614
rect 588542 626378 588778 626614
rect 588222 626058 588458 626294
rect 588542 626058 588778 626294
rect 588222 590378 588458 590614
rect 588542 590378 588778 590614
rect 588222 590058 588458 590294
rect 588542 590058 588778 590294
rect 588222 554378 588458 554614
rect 588542 554378 588778 554614
rect 588222 554058 588458 554294
rect 588542 554058 588778 554294
rect 588222 518378 588458 518614
rect 588542 518378 588778 518614
rect 588222 518058 588458 518294
rect 588542 518058 588778 518294
rect 588222 482378 588458 482614
rect 588542 482378 588778 482614
rect 588222 482058 588458 482294
rect 588542 482058 588778 482294
rect 588222 446378 588458 446614
rect 588542 446378 588778 446614
rect 588222 446058 588458 446294
rect 588542 446058 588778 446294
rect 588222 410378 588458 410614
rect 588542 410378 588778 410614
rect 588222 410058 588458 410294
rect 588542 410058 588778 410294
rect 588222 374378 588458 374614
rect 588542 374378 588778 374614
rect 588222 374058 588458 374294
rect 588542 374058 588778 374294
rect 588222 338378 588458 338614
rect 588542 338378 588778 338614
rect 588222 338058 588458 338294
rect 588542 338058 588778 338294
rect 588222 302378 588458 302614
rect 588542 302378 588778 302614
rect 588222 302058 588458 302294
rect 588542 302058 588778 302294
rect 588222 266378 588458 266614
rect 588542 266378 588778 266614
rect 588222 266058 588458 266294
rect 588542 266058 588778 266294
rect 588222 230378 588458 230614
rect 588542 230378 588778 230614
rect 588222 230058 588458 230294
rect 588542 230058 588778 230294
rect 588222 194378 588458 194614
rect 588542 194378 588778 194614
rect 588222 194058 588458 194294
rect 588542 194058 588778 194294
rect 588222 158378 588458 158614
rect 588542 158378 588778 158614
rect 588222 158058 588458 158294
rect 588542 158058 588778 158294
rect 588222 122378 588458 122614
rect 588542 122378 588778 122614
rect 588222 122058 588458 122294
rect 588542 122058 588778 122294
rect 588222 86378 588458 86614
rect 588542 86378 588778 86614
rect 588222 86058 588458 86294
rect 588542 86058 588778 86294
rect 588222 50378 588458 50614
rect 588542 50378 588778 50614
rect 588222 50058 588458 50294
rect 588542 50058 588778 50294
rect 588222 14378 588458 14614
rect 588542 14378 588778 14614
rect 588222 14058 588458 14294
rect 588542 14058 588778 14294
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 666098 589418 666334
rect 589502 666098 589738 666334
rect 589182 665778 589418 666014
rect 589502 665778 589738 666014
rect 589182 630098 589418 630334
rect 589502 630098 589738 630334
rect 589182 629778 589418 630014
rect 589502 629778 589738 630014
rect 589182 594098 589418 594334
rect 589502 594098 589738 594334
rect 589182 593778 589418 594014
rect 589502 593778 589738 594014
rect 589182 558098 589418 558334
rect 589502 558098 589738 558334
rect 589182 557778 589418 558014
rect 589502 557778 589738 558014
rect 589182 522098 589418 522334
rect 589502 522098 589738 522334
rect 589182 521778 589418 522014
rect 589502 521778 589738 522014
rect 589182 486098 589418 486334
rect 589502 486098 589738 486334
rect 589182 485778 589418 486014
rect 589502 485778 589738 486014
rect 589182 450098 589418 450334
rect 589502 450098 589738 450334
rect 589182 449778 589418 450014
rect 589502 449778 589738 450014
rect 589182 414098 589418 414334
rect 589502 414098 589738 414334
rect 589182 413778 589418 414014
rect 589502 413778 589738 414014
rect 589182 378098 589418 378334
rect 589502 378098 589738 378334
rect 589182 377778 589418 378014
rect 589502 377778 589738 378014
rect 589182 342098 589418 342334
rect 589502 342098 589738 342334
rect 589182 341778 589418 342014
rect 589502 341778 589738 342014
rect 589182 306098 589418 306334
rect 589502 306098 589738 306334
rect 589182 305778 589418 306014
rect 589502 305778 589738 306014
rect 589182 270098 589418 270334
rect 589502 270098 589738 270334
rect 589182 269778 589418 270014
rect 589502 269778 589738 270014
rect 589182 234098 589418 234334
rect 589502 234098 589738 234334
rect 589182 233778 589418 234014
rect 589502 233778 589738 234014
rect 589182 198098 589418 198334
rect 589502 198098 589738 198334
rect 589182 197778 589418 198014
rect 589502 197778 589738 198014
rect 589182 162098 589418 162334
rect 589502 162098 589738 162334
rect 589182 161778 589418 162014
rect 589502 161778 589738 162014
rect 589182 126098 589418 126334
rect 589502 126098 589738 126334
rect 589182 125778 589418 126014
rect 589502 125778 589738 126014
rect 589182 90098 589418 90334
rect 589502 90098 589738 90334
rect 589182 89778 589418 90014
rect 589502 89778 589738 90014
rect 589182 54098 589418 54334
rect 589502 54098 589738 54334
rect 589182 53778 589418 54014
rect 589502 53778 589738 54014
rect 589182 18098 589418 18334
rect 589502 18098 589738 18334
rect 589182 17778 589418 18014
rect 589502 17778 589738 18014
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 669818 590378 670054
rect 590462 669818 590698 670054
rect 590142 669498 590378 669734
rect 590462 669498 590698 669734
rect 590142 633818 590378 634054
rect 590462 633818 590698 634054
rect 590142 633498 590378 633734
rect 590462 633498 590698 633734
rect 590142 597818 590378 598054
rect 590462 597818 590698 598054
rect 590142 597498 590378 597734
rect 590462 597498 590698 597734
rect 590142 561818 590378 562054
rect 590462 561818 590698 562054
rect 590142 561498 590378 561734
rect 590462 561498 590698 561734
rect 590142 525818 590378 526054
rect 590462 525818 590698 526054
rect 590142 525498 590378 525734
rect 590462 525498 590698 525734
rect 590142 489818 590378 490054
rect 590462 489818 590698 490054
rect 590142 489498 590378 489734
rect 590462 489498 590698 489734
rect 590142 453818 590378 454054
rect 590462 453818 590698 454054
rect 590142 453498 590378 453734
rect 590462 453498 590698 453734
rect 590142 417818 590378 418054
rect 590462 417818 590698 418054
rect 590142 417498 590378 417734
rect 590462 417498 590698 417734
rect 590142 381818 590378 382054
rect 590462 381818 590698 382054
rect 590142 381498 590378 381734
rect 590462 381498 590698 381734
rect 590142 345818 590378 346054
rect 590462 345818 590698 346054
rect 590142 345498 590378 345734
rect 590462 345498 590698 345734
rect 590142 309818 590378 310054
rect 590462 309818 590698 310054
rect 590142 309498 590378 309734
rect 590462 309498 590698 309734
rect 590142 273818 590378 274054
rect 590462 273818 590698 274054
rect 590142 273498 590378 273734
rect 590462 273498 590698 273734
rect 590142 237818 590378 238054
rect 590462 237818 590698 238054
rect 590142 237498 590378 237734
rect 590462 237498 590698 237734
rect 590142 201818 590378 202054
rect 590462 201818 590698 202054
rect 590142 201498 590378 201734
rect 590462 201498 590698 201734
rect 590142 165818 590378 166054
rect 590462 165818 590698 166054
rect 590142 165498 590378 165734
rect 590462 165498 590698 165734
rect 590142 129818 590378 130054
rect 590462 129818 590698 130054
rect 590142 129498 590378 129734
rect 590462 129498 590698 129734
rect 590142 93818 590378 94054
rect 590462 93818 590698 94054
rect 590142 93498 590378 93734
rect 590462 93498 590698 93734
rect 590142 57818 590378 58054
rect 590462 57818 590698 58054
rect 590142 57498 590378 57734
rect 590462 57498 590698 57734
rect 590142 21818 590378 22054
rect 590462 21818 590698 22054
rect 590142 21498 590378 21734
rect 590462 21498 590698 21734
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 673538 591338 673774
rect 591422 673538 591658 673774
rect 591102 673218 591338 673454
rect 591422 673218 591658 673454
rect 591102 637538 591338 637774
rect 591422 637538 591658 637774
rect 591102 637218 591338 637454
rect 591422 637218 591658 637454
rect 591102 601538 591338 601774
rect 591422 601538 591658 601774
rect 591102 601218 591338 601454
rect 591422 601218 591658 601454
rect 591102 565538 591338 565774
rect 591422 565538 591658 565774
rect 591102 565218 591338 565454
rect 591422 565218 591658 565454
rect 591102 529538 591338 529774
rect 591422 529538 591658 529774
rect 591102 529218 591338 529454
rect 591422 529218 591658 529454
rect 591102 493538 591338 493774
rect 591422 493538 591658 493774
rect 591102 493218 591338 493454
rect 591422 493218 591658 493454
rect 591102 457538 591338 457774
rect 591422 457538 591658 457774
rect 591102 457218 591338 457454
rect 591422 457218 591658 457454
rect 591102 421538 591338 421774
rect 591422 421538 591658 421774
rect 591102 421218 591338 421454
rect 591422 421218 591658 421454
rect 591102 385538 591338 385774
rect 591422 385538 591658 385774
rect 591102 385218 591338 385454
rect 591422 385218 591658 385454
rect 591102 349538 591338 349774
rect 591422 349538 591658 349774
rect 591102 349218 591338 349454
rect 591422 349218 591658 349454
rect 591102 313538 591338 313774
rect 591422 313538 591658 313774
rect 591102 313218 591338 313454
rect 591422 313218 591658 313454
rect 591102 277538 591338 277774
rect 591422 277538 591658 277774
rect 591102 277218 591338 277454
rect 591422 277218 591658 277454
rect 591102 241538 591338 241774
rect 591422 241538 591658 241774
rect 591102 241218 591338 241454
rect 591422 241218 591658 241454
rect 591102 205538 591338 205774
rect 591422 205538 591658 205774
rect 591102 205218 591338 205454
rect 591422 205218 591658 205454
rect 591102 169538 591338 169774
rect 591422 169538 591658 169774
rect 591102 169218 591338 169454
rect 591422 169218 591658 169454
rect 591102 133538 591338 133774
rect 591422 133538 591658 133774
rect 591102 133218 591338 133454
rect 591422 133218 591658 133454
rect 591102 97538 591338 97774
rect 591422 97538 591658 97774
rect 591102 97218 591338 97454
rect 591422 97218 591658 97454
rect 591102 61538 591338 61774
rect 591422 61538 591658 61774
rect 591102 61218 591338 61454
rect 591422 61218 591658 61454
rect 591102 25538 591338 25774
rect 591422 25538 591658 25774
rect 591102 25218 591338 25454
rect 591422 25218 591658 25454
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 677258 592298 677494
rect 592382 677258 592618 677494
rect 592062 676938 592298 677174
rect 592382 676938 592618 677174
rect 592062 641258 592298 641494
rect 592382 641258 592618 641494
rect 592062 640938 592298 641174
rect 592382 640938 592618 641174
rect 592062 605258 592298 605494
rect 592382 605258 592618 605494
rect 592062 604938 592298 605174
rect 592382 604938 592618 605174
rect 592062 569258 592298 569494
rect 592382 569258 592618 569494
rect 592062 568938 592298 569174
rect 592382 568938 592618 569174
rect 592062 533258 592298 533494
rect 592382 533258 592618 533494
rect 592062 532938 592298 533174
rect 592382 532938 592618 533174
rect 592062 497258 592298 497494
rect 592382 497258 592618 497494
rect 592062 496938 592298 497174
rect 592382 496938 592618 497174
rect 592062 461258 592298 461494
rect 592382 461258 592618 461494
rect 592062 460938 592298 461174
rect 592382 460938 592618 461174
rect 592062 425258 592298 425494
rect 592382 425258 592618 425494
rect 592062 424938 592298 425174
rect 592382 424938 592618 425174
rect 592062 389258 592298 389494
rect 592382 389258 592618 389494
rect 592062 388938 592298 389174
rect 592382 388938 592618 389174
rect 592062 353258 592298 353494
rect 592382 353258 592618 353494
rect 592062 352938 592298 353174
rect 592382 352938 592618 353174
rect 592062 317258 592298 317494
rect 592382 317258 592618 317494
rect 592062 316938 592298 317174
rect 592382 316938 592618 317174
rect 592062 281258 592298 281494
rect 592382 281258 592618 281494
rect 592062 280938 592298 281174
rect 592382 280938 592618 281174
rect 592062 245258 592298 245494
rect 592382 245258 592618 245494
rect 592062 244938 592298 245174
rect 592382 244938 592618 245174
rect 592062 209258 592298 209494
rect 592382 209258 592618 209494
rect 592062 208938 592298 209174
rect 592382 208938 592618 209174
rect 592062 173258 592298 173494
rect 592382 173258 592618 173494
rect 592062 172938 592298 173174
rect 592382 172938 592618 173174
rect 592062 137258 592298 137494
rect 592382 137258 592618 137494
rect 592062 136938 592298 137174
rect 592382 136938 592618 137174
rect 592062 101258 592298 101494
rect 592382 101258 592618 101494
rect 592062 100938 592298 101174
rect 592382 100938 592618 101174
rect 592062 65258 592298 65494
rect 592382 65258 592618 65494
rect 592062 64938 592298 65174
rect 592382 64938 592618 65174
rect 592062 29258 592298 29494
rect 592382 29258 592618 29494
rect 592062 28938 592298 29174
rect 592382 28938 592618 29174
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 12986 707718
rect 13222 707482 13306 707718
rect 13542 707482 48986 707718
rect 49222 707482 49306 707718
rect 49542 707482 84986 707718
rect 85222 707482 85306 707718
rect 85542 707482 120986 707718
rect 121222 707482 121306 707718
rect 121542 707482 156986 707718
rect 157222 707482 157306 707718
rect 157542 707482 192986 707718
rect 193222 707482 193306 707718
rect 193542 707482 228986 707718
rect 229222 707482 229306 707718
rect 229542 707482 264986 707718
rect 265222 707482 265306 707718
rect 265542 707482 300986 707718
rect 301222 707482 301306 707718
rect 301542 707482 336986 707718
rect 337222 707482 337306 707718
rect 337542 707482 372986 707718
rect 373222 707482 373306 707718
rect 373542 707482 408986 707718
rect 409222 707482 409306 707718
rect 409542 707482 444986 707718
rect 445222 707482 445306 707718
rect 445542 707482 480986 707718
rect 481222 707482 481306 707718
rect 481542 707482 516986 707718
rect 517222 707482 517306 707718
rect 517542 707482 552986 707718
rect 553222 707482 553306 707718
rect 553542 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 12986 707398
rect 13222 707162 13306 707398
rect 13542 707162 48986 707398
rect 49222 707162 49306 707398
rect 49542 707162 84986 707398
rect 85222 707162 85306 707398
rect 85542 707162 120986 707398
rect 121222 707162 121306 707398
rect 121542 707162 156986 707398
rect 157222 707162 157306 707398
rect 157542 707162 192986 707398
rect 193222 707162 193306 707398
rect 193542 707162 228986 707398
rect 229222 707162 229306 707398
rect 229542 707162 264986 707398
rect 265222 707162 265306 707398
rect 265542 707162 300986 707398
rect 301222 707162 301306 707398
rect 301542 707162 336986 707398
rect 337222 707162 337306 707398
rect 337542 707162 372986 707398
rect 373222 707162 373306 707398
rect 373542 707162 408986 707398
rect 409222 707162 409306 707398
rect 409542 707162 444986 707398
rect 445222 707162 445306 707398
rect 445542 707162 480986 707398
rect 481222 707162 481306 707398
rect 481542 707162 516986 707398
rect 517222 707162 517306 707398
rect 517542 707162 552986 707398
rect 553222 707162 553306 707398
rect 553542 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 9266 706758
rect 9502 706522 9586 706758
rect 9822 706522 45266 706758
rect 45502 706522 45586 706758
rect 45822 706522 81266 706758
rect 81502 706522 81586 706758
rect 81822 706522 117266 706758
rect 117502 706522 117586 706758
rect 117822 706522 153266 706758
rect 153502 706522 153586 706758
rect 153822 706522 189266 706758
rect 189502 706522 189586 706758
rect 189822 706522 225266 706758
rect 225502 706522 225586 706758
rect 225822 706522 261266 706758
rect 261502 706522 261586 706758
rect 261822 706522 297266 706758
rect 297502 706522 297586 706758
rect 297822 706522 333266 706758
rect 333502 706522 333586 706758
rect 333822 706522 369266 706758
rect 369502 706522 369586 706758
rect 369822 706522 405266 706758
rect 405502 706522 405586 706758
rect 405822 706522 441266 706758
rect 441502 706522 441586 706758
rect 441822 706522 477266 706758
rect 477502 706522 477586 706758
rect 477822 706522 513266 706758
rect 513502 706522 513586 706758
rect 513822 706522 549266 706758
rect 549502 706522 549586 706758
rect 549822 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 9266 706438
rect 9502 706202 9586 706438
rect 9822 706202 45266 706438
rect 45502 706202 45586 706438
rect 45822 706202 81266 706438
rect 81502 706202 81586 706438
rect 81822 706202 117266 706438
rect 117502 706202 117586 706438
rect 117822 706202 153266 706438
rect 153502 706202 153586 706438
rect 153822 706202 189266 706438
rect 189502 706202 189586 706438
rect 189822 706202 225266 706438
rect 225502 706202 225586 706438
rect 225822 706202 261266 706438
rect 261502 706202 261586 706438
rect 261822 706202 297266 706438
rect 297502 706202 297586 706438
rect 297822 706202 333266 706438
rect 333502 706202 333586 706438
rect 333822 706202 369266 706438
rect 369502 706202 369586 706438
rect 369822 706202 405266 706438
rect 405502 706202 405586 706438
rect 405822 706202 441266 706438
rect 441502 706202 441586 706438
rect 441822 706202 477266 706438
rect 477502 706202 477586 706438
rect 477822 706202 513266 706438
rect 513502 706202 513586 706438
rect 513822 706202 549266 706438
rect 549502 706202 549586 706438
rect 549822 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -4854 698614
rect -4618 698378 -4534 698614
rect -4298 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 588222 698614
rect 588458 698378 588542 698614
rect 588778 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -4854 698294
rect -4618 698058 -4534 698294
rect -4298 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 588222 698294
rect 588458 698058 588542 698294
rect 588778 698058 592650 698294
rect -8726 698026 592650 698058
rect -8726 694894 592650 694926
rect -8726 694658 -3894 694894
rect -3658 694658 -3574 694894
rect -3338 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 587262 694894
rect 587498 694658 587582 694894
rect 587818 694658 592650 694894
rect -8726 694574 592650 694658
rect -8726 694338 -3894 694574
rect -3658 694338 -3574 694574
rect -3338 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 587262 694574
rect 587498 694338 587582 694574
rect 587818 694338 592650 694574
rect -8726 694306 592650 694338
rect -8726 691174 592650 691206
rect -8726 690938 -2934 691174
rect -2698 690938 -2614 691174
rect -2378 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 586302 691174
rect 586538 690938 586622 691174
rect 586858 690938 592650 691174
rect -8726 690854 592650 690938
rect -8726 690618 -2934 690854
rect -2698 690618 -2614 690854
rect -2378 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 586302 690854
rect 586538 690618 586622 690854
rect 586858 690618 592650 690854
rect -8726 690586 592650 690618
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 10250 687454
rect 10486 687218 40970 687454
rect 41206 687218 71690 687454
rect 71926 687218 102410 687454
rect 102646 687218 133130 687454
rect 133366 687218 163850 687454
rect 164086 687218 194570 687454
rect 194806 687218 225290 687454
rect 225526 687218 256010 687454
rect 256246 687218 286730 687454
rect 286966 687218 317450 687454
rect 317686 687218 348170 687454
rect 348406 687218 378890 687454
rect 379126 687218 409610 687454
rect 409846 687218 440330 687454
rect 440566 687218 471050 687454
rect 471286 687218 501770 687454
rect 502006 687218 532490 687454
rect 532726 687218 563210 687454
rect 563446 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 10250 687134
rect 10486 686898 40970 687134
rect 41206 686898 71690 687134
rect 71926 686898 102410 687134
rect 102646 686898 133130 687134
rect 133366 686898 163850 687134
rect 164086 686898 194570 687134
rect 194806 686898 225290 687134
rect 225526 686898 256010 687134
rect 256246 686898 286730 687134
rect 286966 686898 317450 687134
rect 317686 686898 348170 687134
rect 348406 686898 378890 687134
rect 379126 686898 409610 687134
rect 409846 686898 440330 687134
rect 440566 686898 471050 687134
rect 471286 686898 501770 687134
rect 502006 686898 532490 687134
rect 532726 686898 563210 687134
rect 563446 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 677494 592650 677526
rect -8726 677258 -8694 677494
rect -8458 677258 -8374 677494
rect -8138 677258 592062 677494
rect 592298 677258 592382 677494
rect 592618 677258 592650 677494
rect -8726 677174 592650 677258
rect -8726 676938 -8694 677174
rect -8458 676938 -8374 677174
rect -8138 676938 592062 677174
rect 592298 676938 592382 677174
rect 592618 676938 592650 677174
rect -8726 676906 592650 676938
rect -8726 673774 592650 673806
rect -8726 673538 -7734 673774
rect -7498 673538 -7414 673774
rect -7178 673538 591102 673774
rect 591338 673538 591422 673774
rect 591658 673538 592650 673774
rect -8726 673454 592650 673538
rect -8726 673218 -7734 673454
rect -7498 673218 -7414 673454
rect -7178 673218 591102 673454
rect 591338 673218 591422 673454
rect 591658 673218 592650 673454
rect -8726 673186 592650 673218
rect -8726 670054 592650 670086
rect -8726 669818 -6774 670054
rect -6538 669818 -6454 670054
rect -6218 669818 590142 670054
rect 590378 669818 590462 670054
rect 590698 669818 592650 670054
rect -8726 669734 592650 669818
rect -8726 669498 -6774 669734
rect -6538 669498 -6454 669734
rect -6218 669498 590142 669734
rect 590378 669498 590462 669734
rect 590698 669498 592650 669734
rect -8726 669466 592650 669498
rect -8726 666334 592650 666366
rect -8726 666098 -5814 666334
rect -5578 666098 -5494 666334
rect -5258 666098 589182 666334
rect 589418 666098 589502 666334
rect 589738 666098 592650 666334
rect -8726 666014 592650 666098
rect -8726 665778 -5814 666014
rect -5578 665778 -5494 666014
rect -5258 665778 589182 666014
rect 589418 665778 589502 666014
rect 589738 665778 592650 666014
rect -8726 665746 592650 665778
rect -8726 662614 592650 662646
rect -8726 662378 -4854 662614
rect -4618 662378 -4534 662614
rect -4298 662378 588222 662614
rect 588458 662378 588542 662614
rect 588778 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -4854 662294
rect -4618 662058 -4534 662294
rect -4298 662058 588222 662294
rect 588458 662058 588542 662294
rect 588778 662058 592650 662294
rect -8726 662026 592650 662058
rect -8726 658894 592650 658926
rect -8726 658658 -3894 658894
rect -3658 658658 -3574 658894
rect -3338 658658 587262 658894
rect 587498 658658 587582 658894
rect 587818 658658 592650 658894
rect -8726 658574 592650 658658
rect -8726 658338 -3894 658574
rect -3658 658338 -3574 658574
rect -3338 658338 587262 658574
rect 587498 658338 587582 658574
rect 587818 658338 592650 658574
rect -8726 658306 592650 658338
rect -8726 655174 592650 655206
rect -8726 654938 -2934 655174
rect -2698 654938 -2614 655174
rect -2378 654938 25610 655174
rect 25846 654938 56330 655174
rect 56566 654938 87050 655174
rect 87286 654938 117770 655174
rect 118006 654938 148490 655174
rect 148726 654938 179210 655174
rect 179446 654938 209930 655174
rect 210166 654938 240650 655174
rect 240886 654938 271370 655174
rect 271606 654938 302090 655174
rect 302326 654938 332810 655174
rect 333046 654938 363530 655174
rect 363766 654938 394250 655174
rect 394486 654938 424970 655174
rect 425206 654938 455690 655174
rect 455926 654938 486410 655174
rect 486646 654938 517130 655174
rect 517366 654938 547850 655174
rect 548086 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 586302 655174
rect 586538 654938 586622 655174
rect 586858 654938 592650 655174
rect -8726 654854 592650 654938
rect -8726 654618 -2934 654854
rect -2698 654618 -2614 654854
rect -2378 654618 25610 654854
rect 25846 654618 56330 654854
rect 56566 654618 87050 654854
rect 87286 654618 117770 654854
rect 118006 654618 148490 654854
rect 148726 654618 179210 654854
rect 179446 654618 209930 654854
rect 210166 654618 240650 654854
rect 240886 654618 271370 654854
rect 271606 654618 302090 654854
rect 302326 654618 332810 654854
rect 333046 654618 363530 654854
rect 363766 654618 394250 654854
rect 394486 654618 424970 654854
rect 425206 654618 455690 654854
rect 455926 654618 486410 654854
rect 486646 654618 517130 654854
rect 517366 654618 547850 654854
rect 548086 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 586302 654854
rect 586538 654618 586622 654854
rect 586858 654618 592650 654854
rect -8726 654586 592650 654618
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 10250 651454
rect 10486 651218 40970 651454
rect 41206 651218 71690 651454
rect 71926 651218 102410 651454
rect 102646 651218 133130 651454
rect 133366 651218 163850 651454
rect 164086 651218 194570 651454
rect 194806 651218 225290 651454
rect 225526 651218 256010 651454
rect 256246 651218 286730 651454
rect 286966 651218 317450 651454
rect 317686 651218 348170 651454
rect 348406 651218 378890 651454
rect 379126 651218 409610 651454
rect 409846 651218 440330 651454
rect 440566 651218 471050 651454
rect 471286 651218 501770 651454
rect 502006 651218 532490 651454
rect 532726 651218 563210 651454
rect 563446 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 10250 651134
rect 10486 650898 40970 651134
rect 41206 650898 71690 651134
rect 71926 650898 102410 651134
rect 102646 650898 133130 651134
rect 133366 650898 163850 651134
rect 164086 650898 194570 651134
rect 194806 650898 225290 651134
rect 225526 650898 256010 651134
rect 256246 650898 286730 651134
rect 286966 650898 317450 651134
rect 317686 650898 348170 651134
rect 348406 650898 378890 651134
rect 379126 650898 409610 651134
rect 409846 650898 440330 651134
rect 440566 650898 471050 651134
rect 471286 650898 501770 651134
rect 502006 650898 532490 651134
rect 532726 650898 563210 651134
rect 563446 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 641494 592650 641526
rect -8726 641258 -8694 641494
rect -8458 641258 -8374 641494
rect -8138 641258 592062 641494
rect 592298 641258 592382 641494
rect 592618 641258 592650 641494
rect -8726 641174 592650 641258
rect -8726 640938 -8694 641174
rect -8458 640938 -8374 641174
rect -8138 640938 592062 641174
rect 592298 640938 592382 641174
rect 592618 640938 592650 641174
rect -8726 640906 592650 640938
rect -8726 637774 592650 637806
rect -8726 637538 -7734 637774
rect -7498 637538 -7414 637774
rect -7178 637538 591102 637774
rect 591338 637538 591422 637774
rect 591658 637538 592650 637774
rect -8726 637454 592650 637538
rect -8726 637218 -7734 637454
rect -7498 637218 -7414 637454
rect -7178 637218 591102 637454
rect 591338 637218 591422 637454
rect 591658 637218 592650 637454
rect -8726 637186 592650 637218
rect -8726 634054 592650 634086
rect -8726 633818 -6774 634054
rect -6538 633818 -6454 634054
rect -6218 633818 590142 634054
rect 590378 633818 590462 634054
rect 590698 633818 592650 634054
rect -8726 633734 592650 633818
rect -8726 633498 -6774 633734
rect -6538 633498 -6454 633734
rect -6218 633498 590142 633734
rect 590378 633498 590462 633734
rect 590698 633498 592650 633734
rect -8726 633466 592650 633498
rect -8726 630334 592650 630366
rect -8726 630098 -5814 630334
rect -5578 630098 -5494 630334
rect -5258 630098 589182 630334
rect 589418 630098 589502 630334
rect 589738 630098 592650 630334
rect -8726 630014 592650 630098
rect -8726 629778 -5814 630014
rect -5578 629778 -5494 630014
rect -5258 629778 589182 630014
rect 589418 629778 589502 630014
rect 589738 629778 592650 630014
rect -8726 629746 592650 629778
rect -8726 626614 592650 626646
rect -8726 626378 -4854 626614
rect -4618 626378 -4534 626614
rect -4298 626378 588222 626614
rect 588458 626378 588542 626614
rect 588778 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -4854 626294
rect -4618 626058 -4534 626294
rect -4298 626058 588222 626294
rect 588458 626058 588542 626294
rect 588778 626058 592650 626294
rect -8726 626026 592650 626058
rect -8726 622894 592650 622926
rect -8726 622658 -3894 622894
rect -3658 622658 -3574 622894
rect -3338 622658 587262 622894
rect 587498 622658 587582 622894
rect 587818 622658 592650 622894
rect -8726 622574 592650 622658
rect -8726 622338 -3894 622574
rect -3658 622338 -3574 622574
rect -3338 622338 587262 622574
rect 587498 622338 587582 622574
rect 587818 622338 592650 622574
rect -8726 622306 592650 622338
rect -8726 619174 592650 619206
rect -8726 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 25610 619174
rect 25846 618938 56330 619174
rect 56566 618938 87050 619174
rect 87286 618938 117770 619174
rect 118006 618938 148490 619174
rect 148726 618938 179210 619174
rect 179446 618938 209930 619174
rect 210166 618938 240650 619174
rect 240886 618938 271370 619174
rect 271606 618938 302090 619174
rect 302326 618938 332810 619174
rect 333046 618938 363530 619174
rect 363766 618938 394250 619174
rect 394486 618938 424970 619174
rect 425206 618938 455690 619174
rect 455926 618938 486410 619174
rect 486646 618938 517130 619174
rect 517366 618938 547850 619174
rect 548086 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 592650 619174
rect -8726 618854 592650 618938
rect -8726 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 25610 618854
rect 25846 618618 56330 618854
rect 56566 618618 87050 618854
rect 87286 618618 117770 618854
rect 118006 618618 148490 618854
rect 148726 618618 179210 618854
rect 179446 618618 209930 618854
rect 210166 618618 240650 618854
rect 240886 618618 271370 618854
rect 271606 618618 302090 618854
rect 302326 618618 332810 618854
rect 333046 618618 363530 618854
rect 363766 618618 394250 618854
rect 394486 618618 424970 618854
rect 425206 618618 455690 618854
rect 455926 618618 486410 618854
rect 486646 618618 517130 618854
rect 517366 618618 547850 618854
rect 548086 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 592650 618854
rect -8726 618586 592650 618618
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 10250 615454
rect 10486 615218 40970 615454
rect 41206 615218 71690 615454
rect 71926 615218 102410 615454
rect 102646 615218 133130 615454
rect 133366 615218 163850 615454
rect 164086 615218 194570 615454
rect 194806 615218 225290 615454
rect 225526 615218 256010 615454
rect 256246 615218 286730 615454
rect 286966 615218 317450 615454
rect 317686 615218 348170 615454
rect 348406 615218 378890 615454
rect 379126 615218 409610 615454
rect 409846 615218 440330 615454
rect 440566 615218 471050 615454
rect 471286 615218 501770 615454
rect 502006 615218 532490 615454
rect 532726 615218 563210 615454
rect 563446 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 10250 615134
rect 10486 614898 40970 615134
rect 41206 614898 71690 615134
rect 71926 614898 102410 615134
rect 102646 614898 133130 615134
rect 133366 614898 163850 615134
rect 164086 614898 194570 615134
rect 194806 614898 225290 615134
rect 225526 614898 256010 615134
rect 256246 614898 286730 615134
rect 286966 614898 317450 615134
rect 317686 614898 348170 615134
rect 348406 614898 378890 615134
rect 379126 614898 409610 615134
rect 409846 614898 440330 615134
rect 440566 614898 471050 615134
rect 471286 614898 501770 615134
rect 502006 614898 532490 615134
rect 532726 614898 563210 615134
rect 563446 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 605494 592650 605526
rect -8726 605258 -8694 605494
rect -8458 605258 -8374 605494
rect -8138 605258 592062 605494
rect 592298 605258 592382 605494
rect 592618 605258 592650 605494
rect -8726 605174 592650 605258
rect -8726 604938 -8694 605174
rect -8458 604938 -8374 605174
rect -8138 604938 592062 605174
rect 592298 604938 592382 605174
rect 592618 604938 592650 605174
rect -8726 604906 592650 604938
rect -8726 601774 592650 601806
rect -8726 601538 -7734 601774
rect -7498 601538 -7414 601774
rect -7178 601538 591102 601774
rect 591338 601538 591422 601774
rect 591658 601538 592650 601774
rect -8726 601454 592650 601538
rect -8726 601218 -7734 601454
rect -7498 601218 -7414 601454
rect -7178 601218 591102 601454
rect 591338 601218 591422 601454
rect 591658 601218 592650 601454
rect -8726 601186 592650 601218
rect -8726 598054 592650 598086
rect -8726 597818 -6774 598054
rect -6538 597818 -6454 598054
rect -6218 597818 590142 598054
rect 590378 597818 590462 598054
rect 590698 597818 592650 598054
rect -8726 597734 592650 597818
rect -8726 597498 -6774 597734
rect -6538 597498 -6454 597734
rect -6218 597498 590142 597734
rect 590378 597498 590462 597734
rect 590698 597498 592650 597734
rect -8726 597466 592650 597498
rect -8726 594334 592650 594366
rect -8726 594098 -5814 594334
rect -5578 594098 -5494 594334
rect -5258 594098 589182 594334
rect 589418 594098 589502 594334
rect 589738 594098 592650 594334
rect -8726 594014 592650 594098
rect -8726 593778 -5814 594014
rect -5578 593778 -5494 594014
rect -5258 593778 589182 594014
rect 589418 593778 589502 594014
rect 589738 593778 592650 594014
rect -8726 593746 592650 593778
rect -8726 590614 592650 590646
rect -8726 590378 -4854 590614
rect -4618 590378 -4534 590614
rect -4298 590378 588222 590614
rect 588458 590378 588542 590614
rect 588778 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -4854 590294
rect -4618 590058 -4534 590294
rect -4298 590058 588222 590294
rect 588458 590058 588542 590294
rect 588778 590058 592650 590294
rect -8726 590026 592650 590058
rect -8726 586894 592650 586926
rect -8726 586658 -3894 586894
rect -3658 586658 -3574 586894
rect -3338 586658 587262 586894
rect 587498 586658 587582 586894
rect 587818 586658 592650 586894
rect -8726 586574 592650 586658
rect -8726 586338 -3894 586574
rect -3658 586338 -3574 586574
rect -3338 586338 587262 586574
rect 587498 586338 587582 586574
rect 587818 586338 592650 586574
rect -8726 586306 592650 586338
rect -8726 583174 592650 583206
rect -8726 582938 -2934 583174
rect -2698 582938 -2614 583174
rect -2378 582938 25610 583174
rect 25846 582938 56330 583174
rect 56566 582938 87050 583174
rect 87286 582938 117770 583174
rect 118006 582938 148490 583174
rect 148726 582938 179210 583174
rect 179446 582938 209930 583174
rect 210166 582938 240650 583174
rect 240886 582938 271370 583174
rect 271606 582938 302090 583174
rect 302326 582938 332810 583174
rect 333046 582938 363530 583174
rect 363766 582938 394250 583174
rect 394486 582938 424970 583174
rect 425206 582938 455690 583174
rect 455926 582938 486410 583174
rect 486646 582938 517130 583174
rect 517366 582938 547850 583174
rect 548086 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 586302 583174
rect 586538 582938 586622 583174
rect 586858 582938 592650 583174
rect -8726 582854 592650 582938
rect -8726 582618 -2934 582854
rect -2698 582618 -2614 582854
rect -2378 582618 25610 582854
rect 25846 582618 56330 582854
rect 56566 582618 87050 582854
rect 87286 582618 117770 582854
rect 118006 582618 148490 582854
rect 148726 582618 179210 582854
rect 179446 582618 209930 582854
rect 210166 582618 240650 582854
rect 240886 582618 271370 582854
rect 271606 582618 302090 582854
rect 302326 582618 332810 582854
rect 333046 582618 363530 582854
rect 363766 582618 394250 582854
rect 394486 582618 424970 582854
rect 425206 582618 455690 582854
rect 455926 582618 486410 582854
rect 486646 582618 517130 582854
rect 517366 582618 547850 582854
rect 548086 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 586302 582854
rect 586538 582618 586622 582854
rect 586858 582618 592650 582854
rect -8726 582586 592650 582618
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 10250 579454
rect 10486 579218 40970 579454
rect 41206 579218 71690 579454
rect 71926 579218 102410 579454
rect 102646 579218 133130 579454
rect 133366 579218 163850 579454
rect 164086 579218 194570 579454
rect 194806 579218 225290 579454
rect 225526 579218 256010 579454
rect 256246 579218 286730 579454
rect 286966 579218 317450 579454
rect 317686 579218 348170 579454
rect 348406 579218 378890 579454
rect 379126 579218 409610 579454
rect 409846 579218 440330 579454
rect 440566 579218 471050 579454
rect 471286 579218 501770 579454
rect 502006 579218 532490 579454
rect 532726 579218 563210 579454
rect 563446 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 10250 579134
rect 10486 578898 40970 579134
rect 41206 578898 71690 579134
rect 71926 578898 102410 579134
rect 102646 578898 133130 579134
rect 133366 578898 163850 579134
rect 164086 578898 194570 579134
rect 194806 578898 225290 579134
rect 225526 578898 256010 579134
rect 256246 578898 286730 579134
rect 286966 578898 317450 579134
rect 317686 578898 348170 579134
rect 348406 578898 378890 579134
rect 379126 578898 409610 579134
rect 409846 578898 440330 579134
rect 440566 578898 471050 579134
rect 471286 578898 501770 579134
rect 502006 578898 532490 579134
rect 532726 578898 563210 579134
rect 563446 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 569494 592650 569526
rect -8726 569258 -8694 569494
rect -8458 569258 -8374 569494
rect -8138 569258 592062 569494
rect 592298 569258 592382 569494
rect 592618 569258 592650 569494
rect -8726 569174 592650 569258
rect -8726 568938 -8694 569174
rect -8458 568938 -8374 569174
rect -8138 568938 592062 569174
rect 592298 568938 592382 569174
rect 592618 568938 592650 569174
rect -8726 568906 592650 568938
rect -8726 565774 592650 565806
rect -8726 565538 -7734 565774
rect -7498 565538 -7414 565774
rect -7178 565538 591102 565774
rect 591338 565538 591422 565774
rect 591658 565538 592650 565774
rect -8726 565454 592650 565538
rect -8726 565218 -7734 565454
rect -7498 565218 -7414 565454
rect -7178 565218 591102 565454
rect 591338 565218 591422 565454
rect 591658 565218 592650 565454
rect -8726 565186 592650 565218
rect -8726 562054 592650 562086
rect -8726 561818 -6774 562054
rect -6538 561818 -6454 562054
rect -6218 561818 590142 562054
rect 590378 561818 590462 562054
rect 590698 561818 592650 562054
rect -8726 561734 592650 561818
rect -8726 561498 -6774 561734
rect -6538 561498 -6454 561734
rect -6218 561498 590142 561734
rect 590378 561498 590462 561734
rect 590698 561498 592650 561734
rect -8726 561466 592650 561498
rect -8726 558334 592650 558366
rect -8726 558098 -5814 558334
rect -5578 558098 -5494 558334
rect -5258 558098 589182 558334
rect 589418 558098 589502 558334
rect 589738 558098 592650 558334
rect -8726 558014 592650 558098
rect -8726 557778 -5814 558014
rect -5578 557778 -5494 558014
rect -5258 557778 589182 558014
rect 589418 557778 589502 558014
rect 589738 557778 592650 558014
rect -8726 557746 592650 557778
rect -8726 554614 592650 554646
rect -8726 554378 -4854 554614
rect -4618 554378 -4534 554614
rect -4298 554378 588222 554614
rect 588458 554378 588542 554614
rect 588778 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -4854 554294
rect -4618 554058 -4534 554294
rect -4298 554058 588222 554294
rect 588458 554058 588542 554294
rect 588778 554058 592650 554294
rect -8726 554026 592650 554058
rect -8726 550894 592650 550926
rect -8726 550658 -3894 550894
rect -3658 550658 -3574 550894
rect -3338 550658 587262 550894
rect 587498 550658 587582 550894
rect 587818 550658 592650 550894
rect -8726 550574 592650 550658
rect -8726 550338 -3894 550574
rect -3658 550338 -3574 550574
rect -3338 550338 587262 550574
rect 587498 550338 587582 550574
rect 587818 550338 592650 550574
rect -8726 550306 592650 550338
rect -8726 547174 592650 547206
rect -8726 546938 -2934 547174
rect -2698 546938 -2614 547174
rect -2378 546938 25610 547174
rect 25846 546938 56330 547174
rect 56566 546938 87050 547174
rect 87286 546938 117770 547174
rect 118006 546938 148490 547174
rect 148726 546938 179210 547174
rect 179446 546938 209930 547174
rect 210166 546938 240650 547174
rect 240886 546938 271370 547174
rect 271606 546938 302090 547174
rect 302326 546938 332810 547174
rect 333046 546938 363530 547174
rect 363766 546938 394250 547174
rect 394486 546938 424970 547174
rect 425206 546938 455690 547174
rect 455926 546938 486410 547174
rect 486646 546938 517130 547174
rect 517366 546938 547850 547174
rect 548086 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 586302 547174
rect 586538 546938 586622 547174
rect 586858 546938 592650 547174
rect -8726 546854 592650 546938
rect -8726 546618 -2934 546854
rect -2698 546618 -2614 546854
rect -2378 546618 25610 546854
rect 25846 546618 56330 546854
rect 56566 546618 87050 546854
rect 87286 546618 117770 546854
rect 118006 546618 148490 546854
rect 148726 546618 179210 546854
rect 179446 546618 209930 546854
rect 210166 546618 240650 546854
rect 240886 546618 271370 546854
rect 271606 546618 302090 546854
rect 302326 546618 332810 546854
rect 333046 546618 363530 546854
rect 363766 546618 394250 546854
rect 394486 546618 424970 546854
rect 425206 546618 455690 546854
rect 455926 546618 486410 546854
rect 486646 546618 517130 546854
rect 517366 546618 547850 546854
rect 548086 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 586302 546854
rect 586538 546618 586622 546854
rect 586858 546618 592650 546854
rect -8726 546586 592650 546618
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 10250 543454
rect 10486 543218 40970 543454
rect 41206 543218 71690 543454
rect 71926 543218 102410 543454
rect 102646 543218 133130 543454
rect 133366 543218 163850 543454
rect 164086 543218 194570 543454
rect 194806 543218 225290 543454
rect 225526 543218 256010 543454
rect 256246 543218 286730 543454
rect 286966 543218 317450 543454
rect 317686 543218 348170 543454
rect 348406 543218 378890 543454
rect 379126 543218 409610 543454
rect 409846 543218 440330 543454
rect 440566 543218 471050 543454
rect 471286 543218 501770 543454
rect 502006 543218 532490 543454
rect 532726 543218 563210 543454
rect 563446 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 10250 543134
rect 10486 542898 40970 543134
rect 41206 542898 71690 543134
rect 71926 542898 102410 543134
rect 102646 542898 133130 543134
rect 133366 542898 163850 543134
rect 164086 542898 194570 543134
rect 194806 542898 225290 543134
rect 225526 542898 256010 543134
rect 256246 542898 286730 543134
rect 286966 542898 317450 543134
rect 317686 542898 348170 543134
rect 348406 542898 378890 543134
rect 379126 542898 409610 543134
rect 409846 542898 440330 543134
rect 440566 542898 471050 543134
rect 471286 542898 501770 543134
rect 502006 542898 532490 543134
rect 532726 542898 563210 543134
rect 563446 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 533494 592650 533526
rect -8726 533258 -8694 533494
rect -8458 533258 -8374 533494
rect -8138 533258 592062 533494
rect 592298 533258 592382 533494
rect 592618 533258 592650 533494
rect -8726 533174 592650 533258
rect -8726 532938 -8694 533174
rect -8458 532938 -8374 533174
rect -8138 532938 592062 533174
rect 592298 532938 592382 533174
rect 592618 532938 592650 533174
rect -8726 532906 592650 532938
rect -8726 529774 592650 529806
rect -8726 529538 -7734 529774
rect -7498 529538 -7414 529774
rect -7178 529538 591102 529774
rect 591338 529538 591422 529774
rect 591658 529538 592650 529774
rect -8726 529454 592650 529538
rect -8726 529218 -7734 529454
rect -7498 529218 -7414 529454
rect -7178 529218 591102 529454
rect 591338 529218 591422 529454
rect 591658 529218 592650 529454
rect -8726 529186 592650 529218
rect -8726 526054 592650 526086
rect -8726 525818 -6774 526054
rect -6538 525818 -6454 526054
rect -6218 525818 590142 526054
rect 590378 525818 590462 526054
rect 590698 525818 592650 526054
rect -8726 525734 592650 525818
rect -8726 525498 -6774 525734
rect -6538 525498 -6454 525734
rect -6218 525498 590142 525734
rect 590378 525498 590462 525734
rect 590698 525498 592650 525734
rect -8726 525466 592650 525498
rect -8726 522334 592650 522366
rect -8726 522098 -5814 522334
rect -5578 522098 -5494 522334
rect -5258 522098 589182 522334
rect 589418 522098 589502 522334
rect 589738 522098 592650 522334
rect -8726 522014 592650 522098
rect -8726 521778 -5814 522014
rect -5578 521778 -5494 522014
rect -5258 521778 589182 522014
rect 589418 521778 589502 522014
rect 589738 521778 592650 522014
rect -8726 521746 592650 521778
rect -8726 518614 592650 518646
rect -8726 518378 -4854 518614
rect -4618 518378 -4534 518614
rect -4298 518378 588222 518614
rect 588458 518378 588542 518614
rect 588778 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -4854 518294
rect -4618 518058 -4534 518294
rect -4298 518058 588222 518294
rect 588458 518058 588542 518294
rect 588778 518058 592650 518294
rect -8726 518026 592650 518058
rect -8726 514894 592650 514926
rect -8726 514658 -3894 514894
rect -3658 514658 -3574 514894
rect -3338 514658 587262 514894
rect 587498 514658 587582 514894
rect 587818 514658 592650 514894
rect -8726 514574 592650 514658
rect -8726 514338 -3894 514574
rect -3658 514338 -3574 514574
rect -3338 514338 587262 514574
rect 587498 514338 587582 514574
rect 587818 514338 592650 514574
rect -8726 514306 592650 514338
rect -8726 511174 592650 511206
rect -8726 510938 -2934 511174
rect -2698 510938 -2614 511174
rect -2378 510938 25610 511174
rect 25846 510938 56330 511174
rect 56566 510938 87050 511174
rect 87286 510938 117770 511174
rect 118006 510938 148490 511174
rect 148726 510938 179210 511174
rect 179446 510938 209930 511174
rect 210166 510938 240650 511174
rect 240886 510938 271370 511174
rect 271606 510938 302090 511174
rect 302326 510938 332810 511174
rect 333046 510938 363530 511174
rect 363766 510938 394250 511174
rect 394486 510938 424970 511174
rect 425206 510938 455690 511174
rect 455926 510938 486410 511174
rect 486646 510938 517130 511174
rect 517366 510938 547850 511174
rect 548086 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 586302 511174
rect 586538 510938 586622 511174
rect 586858 510938 592650 511174
rect -8726 510854 592650 510938
rect -8726 510618 -2934 510854
rect -2698 510618 -2614 510854
rect -2378 510618 25610 510854
rect 25846 510618 56330 510854
rect 56566 510618 87050 510854
rect 87286 510618 117770 510854
rect 118006 510618 148490 510854
rect 148726 510618 179210 510854
rect 179446 510618 209930 510854
rect 210166 510618 240650 510854
rect 240886 510618 271370 510854
rect 271606 510618 302090 510854
rect 302326 510618 332810 510854
rect 333046 510618 363530 510854
rect 363766 510618 394250 510854
rect 394486 510618 424970 510854
rect 425206 510618 455690 510854
rect 455926 510618 486410 510854
rect 486646 510618 517130 510854
rect 517366 510618 547850 510854
rect 548086 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 586302 510854
rect 586538 510618 586622 510854
rect 586858 510618 592650 510854
rect -8726 510586 592650 510618
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 10250 507454
rect 10486 507218 40970 507454
rect 41206 507218 71690 507454
rect 71926 507218 102410 507454
rect 102646 507218 133130 507454
rect 133366 507218 163850 507454
rect 164086 507218 194570 507454
rect 194806 507218 225290 507454
rect 225526 507218 256010 507454
rect 256246 507218 286730 507454
rect 286966 507218 317450 507454
rect 317686 507218 348170 507454
rect 348406 507218 378890 507454
rect 379126 507218 409610 507454
rect 409846 507218 440330 507454
rect 440566 507218 471050 507454
rect 471286 507218 501770 507454
rect 502006 507218 532490 507454
rect 532726 507218 563210 507454
rect 563446 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 10250 507134
rect 10486 506898 40970 507134
rect 41206 506898 71690 507134
rect 71926 506898 102410 507134
rect 102646 506898 133130 507134
rect 133366 506898 163850 507134
rect 164086 506898 194570 507134
rect 194806 506898 225290 507134
rect 225526 506898 256010 507134
rect 256246 506898 286730 507134
rect 286966 506898 317450 507134
rect 317686 506898 348170 507134
rect 348406 506898 378890 507134
rect 379126 506898 409610 507134
rect 409846 506898 440330 507134
rect 440566 506898 471050 507134
rect 471286 506898 501770 507134
rect 502006 506898 532490 507134
rect 532726 506898 563210 507134
rect 563446 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 497494 592650 497526
rect -8726 497258 -8694 497494
rect -8458 497258 -8374 497494
rect -8138 497258 592062 497494
rect 592298 497258 592382 497494
rect 592618 497258 592650 497494
rect -8726 497174 592650 497258
rect -8726 496938 -8694 497174
rect -8458 496938 -8374 497174
rect -8138 496938 592062 497174
rect 592298 496938 592382 497174
rect 592618 496938 592650 497174
rect -8726 496906 592650 496938
rect -8726 493774 592650 493806
rect -8726 493538 -7734 493774
rect -7498 493538 -7414 493774
rect -7178 493538 591102 493774
rect 591338 493538 591422 493774
rect 591658 493538 592650 493774
rect -8726 493454 592650 493538
rect -8726 493218 -7734 493454
rect -7498 493218 -7414 493454
rect -7178 493218 591102 493454
rect 591338 493218 591422 493454
rect 591658 493218 592650 493454
rect -8726 493186 592650 493218
rect -8726 490054 592650 490086
rect -8726 489818 -6774 490054
rect -6538 489818 -6454 490054
rect -6218 489818 590142 490054
rect 590378 489818 590462 490054
rect 590698 489818 592650 490054
rect -8726 489734 592650 489818
rect -8726 489498 -6774 489734
rect -6538 489498 -6454 489734
rect -6218 489498 590142 489734
rect 590378 489498 590462 489734
rect 590698 489498 592650 489734
rect -8726 489466 592650 489498
rect -8726 486334 592650 486366
rect -8726 486098 -5814 486334
rect -5578 486098 -5494 486334
rect -5258 486098 589182 486334
rect 589418 486098 589502 486334
rect 589738 486098 592650 486334
rect -8726 486014 592650 486098
rect -8726 485778 -5814 486014
rect -5578 485778 -5494 486014
rect -5258 485778 589182 486014
rect 589418 485778 589502 486014
rect 589738 485778 592650 486014
rect -8726 485746 592650 485778
rect -8726 482614 592650 482646
rect -8726 482378 -4854 482614
rect -4618 482378 -4534 482614
rect -4298 482378 588222 482614
rect 588458 482378 588542 482614
rect 588778 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -4854 482294
rect -4618 482058 -4534 482294
rect -4298 482058 588222 482294
rect 588458 482058 588542 482294
rect 588778 482058 592650 482294
rect -8726 482026 592650 482058
rect -8726 478894 592650 478926
rect -8726 478658 -3894 478894
rect -3658 478658 -3574 478894
rect -3338 478658 587262 478894
rect 587498 478658 587582 478894
rect 587818 478658 592650 478894
rect -8726 478574 592650 478658
rect -8726 478338 -3894 478574
rect -3658 478338 -3574 478574
rect -3338 478338 587262 478574
rect 587498 478338 587582 478574
rect 587818 478338 592650 478574
rect -8726 478306 592650 478338
rect -8726 475174 592650 475206
rect -8726 474938 -2934 475174
rect -2698 474938 -2614 475174
rect -2378 474938 25610 475174
rect 25846 474938 56330 475174
rect 56566 474938 87050 475174
rect 87286 474938 117770 475174
rect 118006 474938 148490 475174
rect 148726 474938 179210 475174
rect 179446 474938 209930 475174
rect 210166 474938 240650 475174
rect 240886 474938 271370 475174
rect 271606 474938 302090 475174
rect 302326 474938 332810 475174
rect 333046 474938 363530 475174
rect 363766 474938 394250 475174
rect 394486 474938 424970 475174
rect 425206 474938 455690 475174
rect 455926 474938 486410 475174
rect 486646 474938 517130 475174
rect 517366 474938 547850 475174
rect 548086 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 586302 475174
rect 586538 474938 586622 475174
rect 586858 474938 592650 475174
rect -8726 474854 592650 474938
rect -8726 474618 -2934 474854
rect -2698 474618 -2614 474854
rect -2378 474618 25610 474854
rect 25846 474618 56330 474854
rect 56566 474618 87050 474854
rect 87286 474618 117770 474854
rect 118006 474618 148490 474854
rect 148726 474618 179210 474854
rect 179446 474618 209930 474854
rect 210166 474618 240650 474854
rect 240886 474618 271370 474854
rect 271606 474618 302090 474854
rect 302326 474618 332810 474854
rect 333046 474618 363530 474854
rect 363766 474618 394250 474854
rect 394486 474618 424970 474854
rect 425206 474618 455690 474854
rect 455926 474618 486410 474854
rect 486646 474618 517130 474854
rect 517366 474618 547850 474854
rect 548086 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 586302 474854
rect 586538 474618 586622 474854
rect 586858 474618 592650 474854
rect -8726 474586 592650 474618
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 10250 471454
rect 10486 471218 40970 471454
rect 41206 471218 71690 471454
rect 71926 471218 102410 471454
rect 102646 471218 133130 471454
rect 133366 471218 163850 471454
rect 164086 471218 194570 471454
rect 194806 471218 225290 471454
rect 225526 471218 256010 471454
rect 256246 471218 286730 471454
rect 286966 471218 317450 471454
rect 317686 471218 348170 471454
rect 348406 471218 378890 471454
rect 379126 471218 409610 471454
rect 409846 471218 440330 471454
rect 440566 471218 471050 471454
rect 471286 471218 501770 471454
rect 502006 471218 532490 471454
rect 532726 471218 563210 471454
rect 563446 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 10250 471134
rect 10486 470898 40970 471134
rect 41206 470898 71690 471134
rect 71926 470898 102410 471134
rect 102646 470898 133130 471134
rect 133366 470898 163850 471134
rect 164086 470898 194570 471134
rect 194806 470898 225290 471134
rect 225526 470898 256010 471134
rect 256246 470898 286730 471134
rect 286966 470898 317450 471134
rect 317686 470898 348170 471134
rect 348406 470898 378890 471134
rect 379126 470898 409610 471134
rect 409846 470898 440330 471134
rect 440566 470898 471050 471134
rect 471286 470898 501770 471134
rect 502006 470898 532490 471134
rect 532726 470898 563210 471134
rect 563446 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 461494 592650 461526
rect -8726 461258 -8694 461494
rect -8458 461258 -8374 461494
rect -8138 461258 592062 461494
rect 592298 461258 592382 461494
rect 592618 461258 592650 461494
rect -8726 461174 592650 461258
rect -8726 460938 -8694 461174
rect -8458 460938 -8374 461174
rect -8138 460938 592062 461174
rect 592298 460938 592382 461174
rect 592618 460938 592650 461174
rect -8726 460906 592650 460938
rect -8726 457774 592650 457806
rect -8726 457538 -7734 457774
rect -7498 457538 -7414 457774
rect -7178 457538 591102 457774
rect 591338 457538 591422 457774
rect 591658 457538 592650 457774
rect -8726 457454 592650 457538
rect -8726 457218 -7734 457454
rect -7498 457218 -7414 457454
rect -7178 457218 591102 457454
rect 591338 457218 591422 457454
rect 591658 457218 592650 457454
rect -8726 457186 592650 457218
rect -8726 454054 592650 454086
rect -8726 453818 -6774 454054
rect -6538 453818 -6454 454054
rect -6218 453818 590142 454054
rect 590378 453818 590462 454054
rect 590698 453818 592650 454054
rect -8726 453734 592650 453818
rect -8726 453498 -6774 453734
rect -6538 453498 -6454 453734
rect -6218 453498 590142 453734
rect 590378 453498 590462 453734
rect 590698 453498 592650 453734
rect -8726 453466 592650 453498
rect -8726 450334 592650 450366
rect -8726 450098 -5814 450334
rect -5578 450098 -5494 450334
rect -5258 450098 589182 450334
rect 589418 450098 589502 450334
rect 589738 450098 592650 450334
rect -8726 450014 592650 450098
rect -8726 449778 -5814 450014
rect -5578 449778 -5494 450014
rect -5258 449778 589182 450014
rect 589418 449778 589502 450014
rect 589738 449778 592650 450014
rect -8726 449746 592650 449778
rect -8726 446614 592650 446646
rect -8726 446378 -4854 446614
rect -4618 446378 -4534 446614
rect -4298 446378 588222 446614
rect 588458 446378 588542 446614
rect 588778 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -4854 446294
rect -4618 446058 -4534 446294
rect -4298 446058 588222 446294
rect 588458 446058 588542 446294
rect 588778 446058 592650 446294
rect -8726 446026 592650 446058
rect -8726 442894 592650 442926
rect -8726 442658 -3894 442894
rect -3658 442658 -3574 442894
rect -3338 442658 587262 442894
rect 587498 442658 587582 442894
rect 587818 442658 592650 442894
rect -8726 442574 592650 442658
rect -8726 442338 -3894 442574
rect -3658 442338 -3574 442574
rect -3338 442338 587262 442574
rect 587498 442338 587582 442574
rect 587818 442338 592650 442574
rect -8726 442306 592650 442338
rect -8726 439174 592650 439206
rect -8726 438938 -2934 439174
rect -2698 438938 -2614 439174
rect -2378 438938 25610 439174
rect 25846 438938 56330 439174
rect 56566 438938 87050 439174
rect 87286 438938 117770 439174
rect 118006 438938 148490 439174
rect 148726 438938 179210 439174
rect 179446 438938 209930 439174
rect 210166 438938 240650 439174
rect 240886 438938 271370 439174
rect 271606 438938 302090 439174
rect 302326 438938 332810 439174
rect 333046 438938 363530 439174
rect 363766 438938 394250 439174
rect 394486 438938 424970 439174
rect 425206 438938 455690 439174
rect 455926 438938 486410 439174
rect 486646 438938 517130 439174
rect 517366 438938 547850 439174
rect 548086 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 586302 439174
rect 586538 438938 586622 439174
rect 586858 438938 592650 439174
rect -8726 438854 592650 438938
rect -8726 438618 -2934 438854
rect -2698 438618 -2614 438854
rect -2378 438618 25610 438854
rect 25846 438618 56330 438854
rect 56566 438618 87050 438854
rect 87286 438618 117770 438854
rect 118006 438618 148490 438854
rect 148726 438618 179210 438854
rect 179446 438618 209930 438854
rect 210166 438618 240650 438854
rect 240886 438618 271370 438854
rect 271606 438618 302090 438854
rect 302326 438618 332810 438854
rect 333046 438618 363530 438854
rect 363766 438618 394250 438854
rect 394486 438618 424970 438854
rect 425206 438618 455690 438854
rect 455926 438618 486410 438854
rect 486646 438618 517130 438854
rect 517366 438618 547850 438854
rect 548086 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 586302 438854
rect 586538 438618 586622 438854
rect 586858 438618 592650 438854
rect -8726 438586 592650 438618
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 10250 435454
rect 10486 435218 40970 435454
rect 41206 435218 71690 435454
rect 71926 435218 102410 435454
rect 102646 435218 133130 435454
rect 133366 435218 163850 435454
rect 164086 435218 194570 435454
rect 194806 435218 225290 435454
rect 225526 435218 256010 435454
rect 256246 435218 286730 435454
rect 286966 435218 317450 435454
rect 317686 435218 348170 435454
rect 348406 435218 378890 435454
rect 379126 435218 409610 435454
rect 409846 435218 440330 435454
rect 440566 435218 471050 435454
rect 471286 435218 501770 435454
rect 502006 435218 532490 435454
rect 532726 435218 563210 435454
rect 563446 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 10250 435134
rect 10486 434898 40970 435134
rect 41206 434898 71690 435134
rect 71926 434898 102410 435134
rect 102646 434898 133130 435134
rect 133366 434898 163850 435134
rect 164086 434898 194570 435134
rect 194806 434898 225290 435134
rect 225526 434898 256010 435134
rect 256246 434898 286730 435134
rect 286966 434898 317450 435134
rect 317686 434898 348170 435134
rect 348406 434898 378890 435134
rect 379126 434898 409610 435134
rect 409846 434898 440330 435134
rect 440566 434898 471050 435134
rect 471286 434898 501770 435134
rect 502006 434898 532490 435134
rect 532726 434898 563210 435134
rect 563446 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 425494 592650 425526
rect -8726 425258 -8694 425494
rect -8458 425258 -8374 425494
rect -8138 425258 592062 425494
rect 592298 425258 592382 425494
rect 592618 425258 592650 425494
rect -8726 425174 592650 425258
rect -8726 424938 -8694 425174
rect -8458 424938 -8374 425174
rect -8138 424938 592062 425174
rect 592298 424938 592382 425174
rect 592618 424938 592650 425174
rect -8726 424906 592650 424938
rect -8726 421774 592650 421806
rect -8726 421538 -7734 421774
rect -7498 421538 -7414 421774
rect -7178 421538 591102 421774
rect 591338 421538 591422 421774
rect 591658 421538 592650 421774
rect -8726 421454 592650 421538
rect -8726 421218 -7734 421454
rect -7498 421218 -7414 421454
rect -7178 421218 591102 421454
rect 591338 421218 591422 421454
rect 591658 421218 592650 421454
rect -8726 421186 592650 421218
rect -8726 418054 592650 418086
rect -8726 417818 -6774 418054
rect -6538 417818 -6454 418054
rect -6218 417818 590142 418054
rect 590378 417818 590462 418054
rect 590698 417818 592650 418054
rect -8726 417734 592650 417818
rect -8726 417498 -6774 417734
rect -6538 417498 -6454 417734
rect -6218 417498 590142 417734
rect 590378 417498 590462 417734
rect 590698 417498 592650 417734
rect -8726 417466 592650 417498
rect -8726 414334 592650 414366
rect -8726 414098 -5814 414334
rect -5578 414098 -5494 414334
rect -5258 414098 589182 414334
rect 589418 414098 589502 414334
rect 589738 414098 592650 414334
rect -8726 414014 592650 414098
rect -8726 413778 -5814 414014
rect -5578 413778 -5494 414014
rect -5258 413778 589182 414014
rect 589418 413778 589502 414014
rect 589738 413778 592650 414014
rect -8726 413746 592650 413778
rect -8726 410614 592650 410646
rect -8726 410378 -4854 410614
rect -4618 410378 -4534 410614
rect -4298 410378 588222 410614
rect 588458 410378 588542 410614
rect 588778 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -4854 410294
rect -4618 410058 -4534 410294
rect -4298 410058 588222 410294
rect 588458 410058 588542 410294
rect 588778 410058 592650 410294
rect -8726 410026 592650 410058
rect -8726 406894 592650 406926
rect -8726 406658 -3894 406894
rect -3658 406658 -3574 406894
rect -3338 406658 587262 406894
rect 587498 406658 587582 406894
rect 587818 406658 592650 406894
rect -8726 406574 592650 406658
rect -8726 406338 -3894 406574
rect -3658 406338 -3574 406574
rect -3338 406338 587262 406574
rect 587498 406338 587582 406574
rect 587818 406338 592650 406574
rect -8726 406306 592650 406338
rect -8726 403174 592650 403206
rect -8726 402938 -2934 403174
rect -2698 402938 -2614 403174
rect -2378 402938 25610 403174
rect 25846 402938 56330 403174
rect 56566 402938 87050 403174
rect 87286 402938 117770 403174
rect 118006 402938 148490 403174
rect 148726 402938 179210 403174
rect 179446 402938 209930 403174
rect 210166 402938 240650 403174
rect 240886 402938 271370 403174
rect 271606 402938 302090 403174
rect 302326 402938 332810 403174
rect 333046 402938 363530 403174
rect 363766 402938 394250 403174
rect 394486 402938 424970 403174
rect 425206 402938 455690 403174
rect 455926 402938 486410 403174
rect 486646 402938 517130 403174
rect 517366 402938 547850 403174
rect 548086 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 586302 403174
rect 586538 402938 586622 403174
rect 586858 402938 592650 403174
rect -8726 402854 592650 402938
rect -8726 402618 -2934 402854
rect -2698 402618 -2614 402854
rect -2378 402618 25610 402854
rect 25846 402618 56330 402854
rect 56566 402618 87050 402854
rect 87286 402618 117770 402854
rect 118006 402618 148490 402854
rect 148726 402618 179210 402854
rect 179446 402618 209930 402854
rect 210166 402618 240650 402854
rect 240886 402618 271370 402854
rect 271606 402618 302090 402854
rect 302326 402618 332810 402854
rect 333046 402618 363530 402854
rect 363766 402618 394250 402854
rect 394486 402618 424970 402854
rect 425206 402618 455690 402854
rect 455926 402618 486410 402854
rect 486646 402618 517130 402854
rect 517366 402618 547850 402854
rect 548086 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 586302 402854
rect 586538 402618 586622 402854
rect 586858 402618 592650 402854
rect -8726 402586 592650 402618
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 10250 399454
rect 10486 399218 40970 399454
rect 41206 399218 71690 399454
rect 71926 399218 102410 399454
rect 102646 399218 133130 399454
rect 133366 399218 163850 399454
rect 164086 399218 194570 399454
rect 194806 399218 225290 399454
rect 225526 399218 256010 399454
rect 256246 399218 286730 399454
rect 286966 399218 317450 399454
rect 317686 399218 348170 399454
rect 348406 399218 378890 399454
rect 379126 399218 409610 399454
rect 409846 399218 440330 399454
rect 440566 399218 471050 399454
rect 471286 399218 501770 399454
rect 502006 399218 532490 399454
rect 532726 399218 563210 399454
rect 563446 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 10250 399134
rect 10486 398898 40970 399134
rect 41206 398898 71690 399134
rect 71926 398898 102410 399134
rect 102646 398898 133130 399134
rect 133366 398898 163850 399134
rect 164086 398898 194570 399134
rect 194806 398898 225290 399134
rect 225526 398898 256010 399134
rect 256246 398898 286730 399134
rect 286966 398898 317450 399134
rect 317686 398898 348170 399134
rect 348406 398898 378890 399134
rect 379126 398898 409610 399134
rect 409846 398898 440330 399134
rect 440566 398898 471050 399134
rect 471286 398898 501770 399134
rect 502006 398898 532490 399134
rect 532726 398898 563210 399134
rect 563446 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 389494 592650 389526
rect -8726 389258 -8694 389494
rect -8458 389258 -8374 389494
rect -8138 389258 592062 389494
rect 592298 389258 592382 389494
rect 592618 389258 592650 389494
rect -8726 389174 592650 389258
rect -8726 388938 -8694 389174
rect -8458 388938 -8374 389174
rect -8138 388938 592062 389174
rect 592298 388938 592382 389174
rect 592618 388938 592650 389174
rect -8726 388906 592650 388938
rect -8726 385774 592650 385806
rect -8726 385538 -7734 385774
rect -7498 385538 -7414 385774
rect -7178 385538 591102 385774
rect 591338 385538 591422 385774
rect 591658 385538 592650 385774
rect -8726 385454 592650 385538
rect -8726 385218 -7734 385454
rect -7498 385218 -7414 385454
rect -7178 385218 591102 385454
rect 591338 385218 591422 385454
rect 591658 385218 592650 385454
rect -8726 385186 592650 385218
rect -8726 382054 592650 382086
rect -8726 381818 -6774 382054
rect -6538 381818 -6454 382054
rect -6218 381818 590142 382054
rect 590378 381818 590462 382054
rect 590698 381818 592650 382054
rect -8726 381734 592650 381818
rect -8726 381498 -6774 381734
rect -6538 381498 -6454 381734
rect -6218 381498 590142 381734
rect 590378 381498 590462 381734
rect 590698 381498 592650 381734
rect -8726 381466 592650 381498
rect -8726 378334 592650 378366
rect -8726 378098 -5814 378334
rect -5578 378098 -5494 378334
rect -5258 378098 589182 378334
rect 589418 378098 589502 378334
rect 589738 378098 592650 378334
rect -8726 378014 592650 378098
rect -8726 377778 -5814 378014
rect -5578 377778 -5494 378014
rect -5258 377778 589182 378014
rect 589418 377778 589502 378014
rect 589738 377778 592650 378014
rect -8726 377746 592650 377778
rect -8726 374614 592650 374646
rect -8726 374378 -4854 374614
rect -4618 374378 -4534 374614
rect -4298 374378 588222 374614
rect 588458 374378 588542 374614
rect 588778 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -4854 374294
rect -4618 374058 -4534 374294
rect -4298 374058 588222 374294
rect 588458 374058 588542 374294
rect 588778 374058 592650 374294
rect -8726 374026 592650 374058
rect -8726 370894 592650 370926
rect -8726 370658 -3894 370894
rect -3658 370658 -3574 370894
rect -3338 370658 587262 370894
rect 587498 370658 587582 370894
rect 587818 370658 592650 370894
rect -8726 370574 592650 370658
rect -8726 370338 -3894 370574
rect -3658 370338 -3574 370574
rect -3338 370338 587262 370574
rect 587498 370338 587582 370574
rect 587818 370338 592650 370574
rect -8726 370306 592650 370338
rect -8726 367174 592650 367206
rect -8726 366938 -2934 367174
rect -2698 366938 -2614 367174
rect -2378 366938 25610 367174
rect 25846 366938 56330 367174
rect 56566 366938 87050 367174
rect 87286 366938 117770 367174
rect 118006 366938 148490 367174
rect 148726 366938 179210 367174
rect 179446 366938 209930 367174
rect 210166 366938 240650 367174
rect 240886 366938 271370 367174
rect 271606 366938 302090 367174
rect 302326 366938 332810 367174
rect 333046 366938 363530 367174
rect 363766 366938 394250 367174
rect 394486 366938 424970 367174
rect 425206 366938 455690 367174
rect 455926 366938 486410 367174
rect 486646 366938 517130 367174
rect 517366 366938 547850 367174
rect 548086 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 586302 367174
rect 586538 366938 586622 367174
rect 586858 366938 592650 367174
rect -8726 366854 592650 366938
rect -8726 366618 -2934 366854
rect -2698 366618 -2614 366854
rect -2378 366618 25610 366854
rect 25846 366618 56330 366854
rect 56566 366618 87050 366854
rect 87286 366618 117770 366854
rect 118006 366618 148490 366854
rect 148726 366618 179210 366854
rect 179446 366618 209930 366854
rect 210166 366618 240650 366854
rect 240886 366618 271370 366854
rect 271606 366618 302090 366854
rect 302326 366618 332810 366854
rect 333046 366618 363530 366854
rect 363766 366618 394250 366854
rect 394486 366618 424970 366854
rect 425206 366618 455690 366854
rect 455926 366618 486410 366854
rect 486646 366618 517130 366854
rect 517366 366618 547850 366854
rect 548086 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 586302 366854
rect 586538 366618 586622 366854
rect 586858 366618 592650 366854
rect -8726 366586 592650 366618
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 10250 363454
rect 10486 363218 40970 363454
rect 41206 363218 71690 363454
rect 71926 363218 102410 363454
rect 102646 363218 133130 363454
rect 133366 363218 163850 363454
rect 164086 363218 194570 363454
rect 194806 363218 225290 363454
rect 225526 363218 256010 363454
rect 256246 363218 286730 363454
rect 286966 363218 317450 363454
rect 317686 363218 348170 363454
rect 348406 363218 378890 363454
rect 379126 363218 409610 363454
rect 409846 363218 440330 363454
rect 440566 363218 471050 363454
rect 471286 363218 501770 363454
rect 502006 363218 532490 363454
rect 532726 363218 563210 363454
rect 563446 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 10250 363134
rect 10486 362898 40970 363134
rect 41206 362898 71690 363134
rect 71926 362898 102410 363134
rect 102646 362898 133130 363134
rect 133366 362898 163850 363134
rect 164086 362898 194570 363134
rect 194806 362898 225290 363134
rect 225526 362898 256010 363134
rect 256246 362898 286730 363134
rect 286966 362898 317450 363134
rect 317686 362898 348170 363134
rect 348406 362898 378890 363134
rect 379126 362898 409610 363134
rect 409846 362898 440330 363134
rect 440566 362898 471050 363134
rect 471286 362898 501770 363134
rect 502006 362898 532490 363134
rect 532726 362898 563210 363134
rect 563446 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 353494 592650 353526
rect -8726 353258 -8694 353494
rect -8458 353258 -8374 353494
rect -8138 353258 592062 353494
rect 592298 353258 592382 353494
rect 592618 353258 592650 353494
rect -8726 353174 592650 353258
rect -8726 352938 -8694 353174
rect -8458 352938 -8374 353174
rect -8138 352938 592062 353174
rect 592298 352938 592382 353174
rect 592618 352938 592650 353174
rect -8726 352906 592650 352938
rect -8726 349774 592650 349806
rect -8726 349538 -7734 349774
rect -7498 349538 -7414 349774
rect -7178 349538 591102 349774
rect 591338 349538 591422 349774
rect 591658 349538 592650 349774
rect -8726 349454 592650 349538
rect -8726 349218 -7734 349454
rect -7498 349218 -7414 349454
rect -7178 349218 591102 349454
rect 591338 349218 591422 349454
rect 591658 349218 592650 349454
rect -8726 349186 592650 349218
rect -8726 346054 592650 346086
rect -8726 345818 -6774 346054
rect -6538 345818 -6454 346054
rect -6218 345818 590142 346054
rect 590378 345818 590462 346054
rect 590698 345818 592650 346054
rect -8726 345734 592650 345818
rect -8726 345498 -6774 345734
rect -6538 345498 -6454 345734
rect -6218 345498 590142 345734
rect 590378 345498 590462 345734
rect 590698 345498 592650 345734
rect -8726 345466 592650 345498
rect -8726 342334 592650 342366
rect -8726 342098 -5814 342334
rect -5578 342098 -5494 342334
rect -5258 342098 589182 342334
rect 589418 342098 589502 342334
rect 589738 342098 592650 342334
rect -8726 342014 592650 342098
rect -8726 341778 -5814 342014
rect -5578 341778 -5494 342014
rect -5258 341778 589182 342014
rect 589418 341778 589502 342014
rect 589738 341778 592650 342014
rect -8726 341746 592650 341778
rect -8726 338614 592650 338646
rect -8726 338378 -4854 338614
rect -4618 338378 -4534 338614
rect -4298 338378 588222 338614
rect 588458 338378 588542 338614
rect 588778 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -4854 338294
rect -4618 338058 -4534 338294
rect -4298 338058 588222 338294
rect 588458 338058 588542 338294
rect 588778 338058 592650 338294
rect -8726 338026 592650 338058
rect -8726 334894 592650 334926
rect -8726 334658 -3894 334894
rect -3658 334658 -3574 334894
rect -3338 334658 587262 334894
rect 587498 334658 587582 334894
rect 587818 334658 592650 334894
rect -8726 334574 592650 334658
rect -8726 334338 -3894 334574
rect -3658 334338 -3574 334574
rect -3338 334338 587262 334574
rect 587498 334338 587582 334574
rect 587818 334338 592650 334574
rect -8726 334306 592650 334338
rect -8726 331174 592650 331206
rect -8726 330938 -2934 331174
rect -2698 330938 -2614 331174
rect -2378 330938 25610 331174
rect 25846 330938 56330 331174
rect 56566 330938 87050 331174
rect 87286 330938 117770 331174
rect 118006 330938 148490 331174
rect 148726 330938 179210 331174
rect 179446 330938 209930 331174
rect 210166 330938 240650 331174
rect 240886 330938 271370 331174
rect 271606 330938 302090 331174
rect 302326 330938 332810 331174
rect 333046 330938 363530 331174
rect 363766 330938 394250 331174
rect 394486 330938 424970 331174
rect 425206 330938 455690 331174
rect 455926 330938 486410 331174
rect 486646 330938 517130 331174
rect 517366 330938 547850 331174
rect 548086 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 586302 331174
rect 586538 330938 586622 331174
rect 586858 330938 592650 331174
rect -8726 330854 592650 330938
rect -8726 330618 -2934 330854
rect -2698 330618 -2614 330854
rect -2378 330618 25610 330854
rect 25846 330618 56330 330854
rect 56566 330618 87050 330854
rect 87286 330618 117770 330854
rect 118006 330618 148490 330854
rect 148726 330618 179210 330854
rect 179446 330618 209930 330854
rect 210166 330618 240650 330854
rect 240886 330618 271370 330854
rect 271606 330618 302090 330854
rect 302326 330618 332810 330854
rect 333046 330618 363530 330854
rect 363766 330618 394250 330854
rect 394486 330618 424970 330854
rect 425206 330618 455690 330854
rect 455926 330618 486410 330854
rect 486646 330618 517130 330854
rect 517366 330618 547850 330854
rect 548086 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 586302 330854
rect 586538 330618 586622 330854
rect 586858 330618 592650 330854
rect -8726 330586 592650 330618
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 10250 327454
rect 10486 327218 40970 327454
rect 41206 327218 71690 327454
rect 71926 327218 102410 327454
rect 102646 327218 133130 327454
rect 133366 327218 163850 327454
rect 164086 327218 194570 327454
rect 194806 327218 225290 327454
rect 225526 327218 256010 327454
rect 256246 327218 286730 327454
rect 286966 327218 317450 327454
rect 317686 327218 348170 327454
rect 348406 327218 378890 327454
rect 379126 327218 409610 327454
rect 409846 327218 440330 327454
rect 440566 327218 471050 327454
rect 471286 327218 501770 327454
rect 502006 327218 532490 327454
rect 532726 327218 563210 327454
rect 563446 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 10250 327134
rect 10486 326898 40970 327134
rect 41206 326898 71690 327134
rect 71926 326898 102410 327134
rect 102646 326898 133130 327134
rect 133366 326898 163850 327134
rect 164086 326898 194570 327134
rect 194806 326898 225290 327134
rect 225526 326898 256010 327134
rect 256246 326898 286730 327134
rect 286966 326898 317450 327134
rect 317686 326898 348170 327134
rect 348406 326898 378890 327134
rect 379126 326898 409610 327134
rect 409846 326898 440330 327134
rect 440566 326898 471050 327134
rect 471286 326898 501770 327134
rect 502006 326898 532490 327134
rect 532726 326898 563210 327134
rect 563446 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 317494 592650 317526
rect -8726 317258 -8694 317494
rect -8458 317258 -8374 317494
rect -8138 317258 592062 317494
rect 592298 317258 592382 317494
rect 592618 317258 592650 317494
rect -8726 317174 592650 317258
rect -8726 316938 -8694 317174
rect -8458 316938 -8374 317174
rect -8138 316938 592062 317174
rect 592298 316938 592382 317174
rect 592618 316938 592650 317174
rect -8726 316906 592650 316938
rect -8726 313774 592650 313806
rect -8726 313538 -7734 313774
rect -7498 313538 -7414 313774
rect -7178 313538 591102 313774
rect 591338 313538 591422 313774
rect 591658 313538 592650 313774
rect -8726 313454 592650 313538
rect -8726 313218 -7734 313454
rect -7498 313218 -7414 313454
rect -7178 313218 591102 313454
rect 591338 313218 591422 313454
rect 591658 313218 592650 313454
rect -8726 313186 592650 313218
rect -8726 310054 592650 310086
rect -8726 309818 -6774 310054
rect -6538 309818 -6454 310054
rect -6218 309818 590142 310054
rect 590378 309818 590462 310054
rect 590698 309818 592650 310054
rect -8726 309734 592650 309818
rect -8726 309498 -6774 309734
rect -6538 309498 -6454 309734
rect -6218 309498 590142 309734
rect 590378 309498 590462 309734
rect 590698 309498 592650 309734
rect -8726 309466 592650 309498
rect -8726 306334 592650 306366
rect -8726 306098 -5814 306334
rect -5578 306098 -5494 306334
rect -5258 306098 589182 306334
rect 589418 306098 589502 306334
rect 589738 306098 592650 306334
rect -8726 306014 592650 306098
rect -8726 305778 -5814 306014
rect -5578 305778 -5494 306014
rect -5258 305778 589182 306014
rect 589418 305778 589502 306014
rect 589738 305778 592650 306014
rect -8726 305746 592650 305778
rect -8726 302614 592650 302646
rect -8726 302378 -4854 302614
rect -4618 302378 -4534 302614
rect -4298 302378 588222 302614
rect 588458 302378 588542 302614
rect 588778 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -4854 302294
rect -4618 302058 -4534 302294
rect -4298 302058 588222 302294
rect 588458 302058 588542 302294
rect 588778 302058 592650 302294
rect -8726 302026 592650 302058
rect -8726 298894 592650 298926
rect -8726 298658 -3894 298894
rect -3658 298658 -3574 298894
rect -3338 298658 587262 298894
rect 587498 298658 587582 298894
rect 587818 298658 592650 298894
rect -8726 298574 592650 298658
rect -8726 298338 -3894 298574
rect -3658 298338 -3574 298574
rect -3338 298338 587262 298574
rect 587498 298338 587582 298574
rect 587818 298338 592650 298574
rect -8726 298306 592650 298338
rect -8726 295174 592650 295206
rect -8726 294938 -2934 295174
rect -2698 294938 -2614 295174
rect -2378 294938 25610 295174
rect 25846 294938 56330 295174
rect 56566 294938 87050 295174
rect 87286 294938 117770 295174
rect 118006 294938 148490 295174
rect 148726 294938 179210 295174
rect 179446 294938 209930 295174
rect 210166 294938 240650 295174
rect 240886 294938 271370 295174
rect 271606 294938 302090 295174
rect 302326 294938 332810 295174
rect 333046 294938 363530 295174
rect 363766 294938 394250 295174
rect 394486 294938 424970 295174
rect 425206 294938 455690 295174
rect 455926 294938 486410 295174
rect 486646 294938 517130 295174
rect 517366 294938 547850 295174
rect 548086 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 586302 295174
rect 586538 294938 586622 295174
rect 586858 294938 592650 295174
rect -8726 294854 592650 294938
rect -8726 294618 -2934 294854
rect -2698 294618 -2614 294854
rect -2378 294618 25610 294854
rect 25846 294618 56330 294854
rect 56566 294618 87050 294854
rect 87286 294618 117770 294854
rect 118006 294618 148490 294854
rect 148726 294618 179210 294854
rect 179446 294618 209930 294854
rect 210166 294618 240650 294854
rect 240886 294618 271370 294854
rect 271606 294618 302090 294854
rect 302326 294618 332810 294854
rect 333046 294618 363530 294854
rect 363766 294618 394250 294854
rect 394486 294618 424970 294854
rect 425206 294618 455690 294854
rect 455926 294618 486410 294854
rect 486646 294618 517130 294854
rect 517366 294618 547850 294854
rect 548086 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 586302 294854
rect 586538 294618 586622 294854
rect 586858 294618 592650 294854
rect -8726 294586 592650 294618
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 10250 291454
rect 10486 291218 40970 291454
rect 41206 291218 71690 291454
rect 71926 291218 102410 291454
rect 102646 291218 133130 291454
rect 133366 291218 163850 291454
rect 164086 291218 194570 291454
rect 194806 291218 225290 291454
rect 225526 291218 256010 291454
rect 256246 291218 286730 291454
rect 286966 291218 317450 291454
rect 317686 291218 348170 291454
rect 348406 291218 378890 291454
rect 379126 291218 409610 291454
rect 409846 291218 440330 291454
rect 440566 291218 471050 291454
rect 471286 291218 501770 291454
rect 502006 291218 532490 291454
rect 532726 291218 563210 291454
rect 563446 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 10250 291134
rect 10486 290898 40970 291134
rect 41206 290898 71690 291134
rect 71926 290898 102410 291134
rect 102646 290898 133130 291134
rect 133366 290898 163850 291134
rect 164086 290898 194570 291134
rect 194806 290898 225290 291134
rect 225526 290898 256010 291134
rect 256246 290898 286730 291134
rect 286966 290898 317450 291134
rect 317686 290898 348170 291134
rect 348406 290898 378890 291134
rect 379126 290898 409610 291134
rect 409846 290898 440330 291134
rect 440566 290898 471050 291134
rect 471286 290898 501770 291134
rect 502006 290898 532490 291134
rect 532726 290898 563210 291134
rect 563446 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 281494 592650 281526
rect -8726 281258 -8694 281494
rect -8458 281258 -8374 281494
rect -8138 281258 592062 281494
rect 592298 281258 592382 281494
rect 592618 281258 592650 281494
rect -8726 281174 592650 281258
rect -8726 280938 -8694 281174
rect -8458 280938 -8374 281174
rect -8138 280938 592062 281174
rect 592298 280938 592382 281174
rect 592618 280938 592650 281174
rect -8726 280906 592650 280938
rect -8726 277774 592650 277806
rect -8726 277538 -7734 277774
rect -7498 277538 -7414 277774
rect -7178 277538 591102 277774
rect 591338 277538 591422 277774
rect 591658 277538 592650 277774
rect -8726 277454 592650 277538
rect -8726 277218 -7734 277454
rect -7498 277218 -7414 277454
rect -7178 277218 591102 277454
rect 591338 277218 591422 277454
rect 591658 277218 592650 277454
rect -8726 277186 592650 277218
rect -8726 274054 592650 274086
rect -8726 273818 -6774 274054
rect -6538 273818 -6454 274054
rect -6218 273818 590142 274054
rect 590378 273818 590462 274054
rect 590698 273818 592650 274054
rect -8726 273734 592650 273818
rect -8726 273498 -6774 273734
rect -6538 273498 -6454 273734
rect -6218 273498 590142 273734
rect 590378 273498 590462 273734
rect 590698 273498 592650 273734
rect -8726 273466 592650 273498
rect -8726 270334 592650 270366
rect -8726 270098 -5814 270334
rect -5578 270098 -5494 270334
rect -5258 270098 589182 270334
rect 589418 270098 589502 270334
rect 589738 270098 592650 270334
rect -8726 270014 592650 270098
rect -8726 269778 -5814 270014
rect -5578 269778 -5494 270014
rect -5258 269778 589182 270014
rect 589418 269778 589502 270014
rect 589738 269778 592650 270014
rect -8726 269746 592650 269778
rect -8726 266614 592650 266646
rect -8726 266378 -4854 266614
rect -4618 266378 -4534 266614
rect -4298 266378 588222 266614
rect 588458 266378 588542 266614
rect 588778 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -4854 266294
rect -4618 266058 -4534 266294
rect -4298 266058 588222 266294
rect 588458 266058 588542 266294
rect 588778 266058 592650 266294
rect -8726 266026 592650 266058
rect -8726 262894 592650 262926
rect -8726 262658 -3894 262894
rect -3658 262658 -3574 262894
rect -3338 262658 587262 262894
rect 587498 262658 587582 262894
rect 587818 262658 592650 262894
rect -8726 262574 592650 262658
rect -8726 262338 -3894 262574
rect -3658 262338 -3574 262574
rect -3338 262338 587262 262574
rect 587498 262338 587582 262574
rect 587818 262338 592650 262574
rect -8726 262306 592650 262338
rect -8726 259174 592650 259206
rect -8726 258938 -2934 259174
rect -2698 258938 -2614 259174
rect -2378 258938 25610 259174
rect 25846 258938 56330 259174
rect 56566 258938 87050 259174
rect 87286 258938 117770 259174
rect 118006 258938 148490 259174
rect 148726 258938 179210 259174
rect 179446 258938 209930 259174
rect 210166 258938 240650 259174
rect 240886 258938 271370 259174
rect 271606 258938 302090 259174
rect 302326 258938 332810 259174
rect 333046 258938 363530 259174
rect 363766 258938 394250 259174
rect 394486 258938 424970 259174
rect 425206 258938 455690 259174
rect 455926 258938 486410 259174
rect 486646 258938 517130 259174
rect 517366 258938 547850 259174
rect 548086 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 586302 259174
rect 586538 258938 586622 259174
rect 586858 258938 592650 259174
rect -8726 258854 592650 258938
rect -8726 258618 -2934 258854
rect -2698 258618 -2614 258854
rect -2378 258618 25610 258854
rect 25846 258618 56330 258854
rect 56566 258618 87050 258854
rect 87286 258618 117770 258854
rect 118006 258618 148490 258854
rect 148726 258618 179210 258854
rect 179446 258618 209930 258854
rect 210166 258618 240650 258854
rect 240886 258618 271370 258854
rect 271606 258618 302090 258854
rect 302326 258618 332810 258854
rect 333046 258618 363530 258854
rect 363766 258618 394250 258854
rect 394486 258618 424970 258854
rect 425206 258618 455690 258854
rect 455926 258618 486410 258854
rect 486646 258618 517130 258854
rect 517366 258618 547850 258854
rect 548086 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 586302 258854
rect 586538 258618 586622 258854
rect 586858 258618 592650 258854
rect -8726 258586 592650 258618
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 10250 255454
rect 10486 255218 40970 255454
rect 41206 255218 71690 255454
rect 71926 255218 102410 255454
rect 102646 255218 133130 255454
rect 133366 255218 163850 255454
rect 164086 255218 194570 255454
rect 194806 255218 225290 255454
rect 225526 255218 256010 255454
rect 256246 255218 286730 255454
rect 286966 255218 317450 255454
rect 317686 255218 348170 255454
rect 348406 255218 378890 255454
rect 379126 255218 409610 255454
rect 409846 255218 440330 255454
rect 440566 255218 471050 255454
rect 471286 255218 501770 255454
rect 502006 255218 532490 255454
rect 532726 255218 563210 255454
rect 563446 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 10250 255134
rect 10486 254898 40970 255134
rect 41206 254898 71690 255134
rect 71926 254898 102410 255134
rect 102646 254898 133130 255134
rect 133366 254898 163850 255134
rect 164086 254898 194570 255134
rect 194806 254898 225290 255134
rect 225526 254898 256010 255134
rect 256246 254898 286730 255134
rect 286966 254898 317450 255134
rect 317686 254898 348170 255134
rect 348406 254898 378890 255134
rect 379126 254898 409610 255134
rect 409846 254898 440330 255134
rect 440566 254898 471050 255134
rect 471286 254898 501770 255134
rect 502006 254898 532490 255134
rect 532726 254898 563210 255134
rect 563446 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 245494 592650 245526
rect -8726 245258 -8694 245494
rect -8458 245258 -8374 245494
rect -8138 245258 592062 245494
rect 592298 245258 592382 245494
rect 592618 245258 592650 245494
rect -8726 245174 592650 245258
rect -8726 244938 -8694 245174
rect -8458 244938 -8374 245174
rect -8138 244938 592062 245174
rect 592298 244938 592382 245174
rect 592618 244938 592650 245174
rect -8726 244906 592650 244938
rect -8726 241774 592650 241806
rect -8726 241538 -7734 241774
rect -7498 241538 -7414 241774
rect -7178 241538 591102 241774
rect 591338 241538 591422 241774
rect 591658 241538 592650 241774
rect -8726 241454 592650 241538
rect -8726 241218 -7734 241454
rect -7498 241218 -7414 241454
rect -7178 241218 591102 241454
rect 591338 241218 591422 241454
rect 591658 241218 592650 241454
rect -8726 241186 592650 241218
rect -8726 238054 592650 238086
rect -8726 237818 -6774 238054
rect -6538 237818 -6454 238054
rect -6218 237818 590142 238054
rect 590378 237818 590462 238054
rect 590698 237818 592650 238054
rect -8726 237734 592650 237818
rect -8726 237498 -6774 237734
rect -6538 237498 -6454 237734
rect -6218 237498 590142 237734
rect 590378 237498 590462 237734
rect 590698 237498 592650 237734
rect -8726 237466 592650 237498
rect -8726 234334 592650 234366
rect -8726 234098 -5814 234334
rect -5578 234098 -5494 234334
rect -5258 234098 589182 234334
rect 589418 234098 589502 234334
rect 589738 234098 592650 234334
rect -8726 234014 592650 234098
rect -8726 233778 -5814 234014
rect -5578 233778 -5494 234014
rect -5258 233778 589182 234014
rect 589418 233778 589502 234014
rect 589738 233778 592650 234014
rect -8726 233746 592650 233778
rect -8726 230614 592650 230646
rect -8726 230378 -4854 230614
rect -4618 230378 -4534 230614
rect -4298 230378 588222 230614
rect 588458 230378 588542 230614
rect 588778 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -4854 230294
rect -4618 230058 -4534 230294
rect -4298 230058 588222 230294
rect 588458 230058 588542 230294
rect 588778 230058 592650 230294
rect -8726 230026 592650 230058
rect -8726 226894 592650 226926
rect -8726 226658 -3894 226894
rect -3658 226658 -3574 226894
rect -3338 226658 587262 226894
rect 587498 226658 587582 226894
rect 587818 226658 592650 226894
rect -8726 226574 592650 226658
rect -8726 226338 -3894 226574
rect -3658 226338 -3574 226574
rect -3338 226338 587262 226574
rect 587498 226338 587582 226574
rect 587818 226338 592650 226574
rect -8726 226306 592650 226338
rect -8726 223174 592650 223206
rect -8726 222938 -2934 223174
rect -2698 222938 -2614 223174
rect -2378 222938 25610 223174
rect 25846 222938 56330 223174
rect 56566 222938 87050 223174
rect 87286 222938 117770 223174
rect 118006 222938 148490 223174
rect 148726 222938 179210 223174
rect 179446 222938 209930 223174
rect 210166 222938 240650 223174
rect 240886 222938 271370 223174
rect 271606 222938 302090 223174
rect 302326 222938 332810 223174
rect 333046 222938 363530 223174
rect 363766 222938 394250 223174
rect 394486 222938 424970 223174
rect 425206 222938 455690 223174
rect 455926 222938 486410 223174
rect 486646 222938 517130 223174
rect 517366 222938 547850 223174
rect 548086 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 586302 223174
rect 586538 222938 586622 223174
rect 586858 222938 592650 223174
rect -8726 222854 592650 222938
rect -8726 222618 -2934 222854
rect -2698 222618 -2614 222854
rect -2378 222618 25610 222854
rect 25846 222618 56330 222854
rect 56566 222618 87050 222854
rect 87286 222618 117770 222854
rect 118006 222618 148490 222854
rect 148726 222618 179210 222854
rect 179446 222618 209930 222854
rect 210166 222618 240650 222854
rect 240886 222618 271370 222854
rect 271606 222618 302090 222854
rect 302326 222618 332810 222854
rect 333046 222618 363530 222854
rect 363766 222618 394250 222854
rect 394486 222618 424970 222854
rect 425206 222618 455690 222854
rect 455926 222618 486410 222854
rect 486646 222618 517130 222854
rect 517366 222618 547850 222854
rect 548086 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 586302 222854
rect 586538 222618 586622 222854
rect 586858 222618 592650 222854
rect -8726 222586 592650 222618
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 10250 219454
rect 10486 219218 40970 219454
rect 41206 219218 71690 219454
rect 71926 219218 102410 219454
rect 102646 219218 133130 219454
rect 133366 219218 163850 219454
rect 164086 219218 194570 219454
rect 194806 219218 225290 219454
rect 225526 219218 256010 219454
rect 256246 219218 286730 219454
rect 286966 219218 317450 219454
rect 317686 219218 348170 219454
rect 348406 219218 378890 219454
rect 379126 219218 409610 219454
rect 409846 219218 440330 219454
rect 440566 219218 471050 219454
rect 471286 219218 501770 219454
rect 502006 219218 532490 219454
rect 532726 219218 563210 219454
rect 563446 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 10250 219134
rect 10486 218898 40970 219134
rect 41206 218898 71690 219134
rect 71926 218898 102410 219134
rect 102646 218898 133130 219134
rect 133366 218898 163850 219134
rect 164086 218898 194570 219134
rect 194806 218898 225290 219134
rect 225526 218898 256010 219134
rect 256246 218898 286730 219134
rect 286966 218898 317450 219134
rect 317686 218898 348170 219134
rect 348406 218898 378890 219134
rect 379126 218898 409610 219134
rect 409846 218898 440330 219134
rect 440566 218898 471050 219134
rect 471286 218898 501770 219134
rect 502006 218898 532490 219134
rect 532726 218898 563210 219134
rect 563446 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 209494 592650 209526
rect -8726 209258 -8694 209494
rect -8458 209258 -8374 209494
rect -8138 209258 592062 209494
rect 592298 209258 592382 209494
rect 592618 209258 592650 209494
rect -8726 209174 592650 209258
rect -8726 208938 -8694 209174
rect -8458 208938 -8374 209174
rect -8138 208938 592062 209174
rect 592298 208938 592382 209174
rect 592618 208938 592650 209174
rect -8726 208906 592650 208938
rect -8726 205774 592650 205806
rect -8726 205538 -7734 205774
rect -7498 205538 -7414 205774
rect -7178 205538 591102 205774
rect 591338 205538 591422 205774
rect 591658 205538 592650 205774
rect -8726 205454 592650 205538
rect -8726 205218 -7734 205454
rect -7498 205218 -7414 205454
rect -7178 205218 591102 205454
rect 591338 205218 591422 205454
rect 591658 205218 592650 205454
rect -8726 205186 592650 205218
rect -8726 202054 592650 202086
rect -8726 201818 -6774 202054
rect -6538 201818 -6454 202054
rect -6218 201818 590142 202054
rect 590378 201818 590462 202054
rect 590698 201818 592650 202054
rect -8726 201734 592650 201818
rect -8726 201498 -6774 201734
rect -6538 201498 -6454 201734
rect -6218 201498 590142 201734
rect 590378 201498 590462 201734
rect 590698 201498 592650 201734
rect -8726 201466 592650 201498
rect -8726 198334 592650 198366
rect -8726 198098 -5814 198334
rect -5578 198098 -5494 198334
rect -5258 198098 589182 198334
rect 589418 198098 589502 198334
rect 589738 198098 592650 198334
rect -8726 198014 592650 198098
rect -8726 197778 -5814 198014
rect -5578 197778 -5494 198014
rect -5258 197778 589182 198014
rect 589418 197778 589502 198014
rect 589738 197778 592650 198014
rect -8726 197746 592650 197778
rect -8726 194614 592650 194646
rect -8726 194378 -4854 194614
rect -4618 194378 -4534 194614
rect -4298 194378 588222 194614
rect 588458 194378 588542 194614
rect 588778 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -4854 194294
rect -4618 194058 -4534 194294
rect -4298 194058 588222 194294
rect 588458 194058 588542 194294
rect 588778 194058 592650 194294
rect -8726 194026 592650 194058
rect -8726 190894 592650 190926
rect -8726 190658 -3894 190894
rect -3658 190658 -3574 190894
rect -3338 190658 587262 190894
rect 587498 190658 587582 190894
rect 587818 190658 592650 190894
rect -8726 190574 592650 190658
rect -8726 190338 -3894 190574
rect -3658 190338 -3574 190574
rect -3338 190338 587262 190574
rect 587498 190338 587582 190574
rect 587818 190338 592650 190574
rect -8726 190306 592650 190338
rect -8726 187174 592650 187206
rect -8726 186938 -2934 187174
rect -2698 186938 -2614 187174
rect -2378 186938 25610 187174
rect 25846 186938 56330 187174
rect 56566 186938 87050 187174
rect 87286 186938 117770 187174
rect 118006 186938 148490 187174
rect 148726 186938 179210 187174
rect 179446 186938 209930 187174
rect 210166 186938 240650 187174
rect 240886 186938 271370 187174
rect 271606 186938 302090 187174
rect 302326 186938 332810 187174
rect 333046 186938 363530 187174
rect 363766 186938 394250 187174
rect 394486 186938 424970 187174
rect 425206 186938 455690 187174
rect 455926 186938 486410 187174
rect 486646 186938 517130 187174
rect 517366 186938 547850 187174
rect 548086 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 586302 187174
rect 586538 186938 586622 187174
rect 586858 186938 592650 187174
rect -8726 186854 592650 186938
rect -8726 186618 -2934 186854
rect -2698 186618 -2614 186854
rect -2378 186618 25610 186854
rect 25846 186618 56330 186854
rect 56566 186618 87050 186854
rect 87286 186618 117770 186854
rect 118006 186618 148490 186854
rect 148726 186618 179210 186854
rect 179446 186618 209930 186854
rect 210166 186618 240650 186854
rect 240886 186618 271370 186854
rect 271606 186618 302090 186854
rect 302326 186618 332810 186854
rect 333046 186618 363530 186854
rect 363766 186618 394250 186854
rect 394486 186618 424970 186854
rect 425206 186618 455690 186854
rect 455926 186618 486410 186854
rect 486646 186618 517130 186854
rect 517366 186618 547850 186854
rect 548086 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 586302 186854
rect 586538 186618 586622 186854
rect 586858 186618 592650 186854
rect -8726 186586 592650 186618
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 10250 183454
rect 10486 183218 40970 183454
rect 41206 183218 71690 183454
rect 71926 183218 102410 183454
rect 102646 183218 133130 183454
rect 133366 183218 163850 183454
rect 164086 183218 194570 183454
rect 194806 183218 225290 183454
rect 225526 183218 256010 183454
rect 256246 183218 286730 183454
rect 286966 183218 317450 183454
rect 317686 183218 348170 183454
rect 348406 183218 378890 183454
rect 379126 183218 409610 183454
rect 409846 183218 440330 183454
rect 440566 183218 471050 183454
rect 471286 183218 501770 183454
rect 502006 183218 532490 183454
rect 532726 183218 563210 183454
rect 563446 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 10250 183134
rect 10486 182898 40970 183134
rect 41206 182898 71690 183134
rect 71926 182898 102410 183134
rect 102646 182898 133130 183134
rect 133366 182898 163850 183134
rect 164086 182898 194570 183134
rect 194806 182898 225290 183134
rect 225526 182898 256010 183134
rect 256246 182898 286730 183134
rect 286966 182898 317450 183134
rect 317686 182898 348170 183134
rect 348406 182898 378890 183134
rect 379126 182898 409610 183134
rect 409846 182898 440330 183134
rect 440566 182898 471050 183134
rect 471286 182898 501770 183134
rect 502006 182898 532490 183134
rect 532726 182898 563210 183134
rect 563446 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 173494 592650 173526
rect -8726 173258 -8694 173494
rect -8458 173258 -8374 173494
rect -8138 173258 592062 173494
rect 592298 173258 592382 173494
rect 592618 173258 592650 173494
rect -8726 173174 592650 173258
rect -8726 172938 -8694 173174
rect -8458 172938 -8374 173174
rect -8138 172938 592062 173174
rect 592298 172938 592382 173174
rect 592618 172938 592650 173174
rect -8726 172906 592650 172938
rect -8726 169774 592650 169806
rect -8726 169538 -7734 169774
rect -7498 169538 -7414 169774
rect -7178 169538 591102 169774
rect 591338 169538 591422 169774
rect 591658 169538 592650 169774
rect -8726 169454 592650 169538
rect -8726 169218 -7734 169454
rect -7498 169218 -7414 169454
rect -7178 169218 591102 169454
rect 591338 169218 591422 169454
rect 591658 169218 592650 169454
rect -8726 169186 592650 169218
rect -8726 166054 592650 166086
rect -8726 165818 -6774 166054
rect -6538 165818 -6454 166054
rect -6218 165818 590142 166054
rect 590378 165818 590462 166054
rect 590698 165818 592650 166054
rect -8726 165734 592650 165818
rect -8726 165498 -6774 165734
rect -6538 165498 -6454 165734
rect -6218 165498 590142 165734
rect 590378 165498 590462 165734
rect 590698 165498 592650 165734
rect -8726 165466 592650 165498
rect -8726 162334 592650 162366
rect -8726 162098 -5814 162334
rect -5578 162098 -5494 162334
rect -5258 162098 589182 162334
rect 589418 162098 589502 162334
rect 589738 162098 592650 162334
rect -8726 162014 592650 162098
rect -8726 161778 -5814 162014
rect -5578 161778 -5494 162014
rect -5258 161778 589182 162014
rect 589418 161778 589502 162014
rect 589738 161778 592650 162014
rect -8726 161746 592650 161778
rect -8726 158614 592650 158646
rect -8726 158378 -4854 158614
rect -4618 158378 -4534 158614
rect -4298 158378 588222 158614
rect 588458 158378 588542 158614
rect 588778 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -4854 158294
rect -4618 158058 -4534 158294
rect -4298 158058 588222 158294
rect 588458 158058 588542 158294
rect 588778 158058 592650 158294
rect -8726 158026 592650 158058
rect -8726 154894 592650 154926
rect -8726 154658 -3894 154894
rect -3658 154658 -3574 154894
rect -3338 154658 587262 154894
rect 587498 154658 587582 154894
rect 587818 154658 592650 154894
rect -8726 154574 592650 154658
rect -8726 154338 -3894 154574
rect -3658 154338 -3574 154574
rect -3338 154338 587262 154574
rect 587498 154338 587582 154574
rect 587818 154338 592650 154574
rect -8726 154306 592650 154338
rect -8726 151174 592650 151206
rect -8726 150938 -2934 151174
rect -2698 150938 -2614 151174
rect -2378 150938 25610 151174
rect 25846 150938 56330 151174
rect 56566 150938 87050 151174
rect 87286 150938 117770 151174
rect 118006 150938 148490 151174
rect 148726 150938 179210 151174
rect 179446 150938 209930 151174
rect 210166 150938 240650 151174
rect 240886 150938 271370 151174
rect 271606 150938 302090 151174
rect 302326 150938 332810 151174
rect 333046 150938 363530 151174
rect 363766 150938 394250 151174
rect 394486 150938 424970 151174
rect 425206 150938 455690 151174
rect 455926 150938 486410 151174
rect 486646 150938 517130 151174
rect 517366 150938 547850 151174
rect 548086 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 586302 151174
rect 586538 150938 586622 151174
rect 586858 150938 592650 151174
rect -8726 150854 592650 150938
rect -8726 150618 -2934 150854
rect -2698 150618 -2614 150854
rect -2378 150618 25610 150854
rect 25846 150618 56330 150854
rect 56566 150618 87050 150854
rect 87286 150618 117770 150854
rect 118006 150618 148490 150854
rect 148726 150618 179210 150854
rect 179446 150618 209930 150854
rect 210166 150618 240650 150854
rect 240886 150618 271370 150854
rect 271606 150618 302090 150854
rect 302326 150618 332810 150854
rect 333046 150618 363530 150854
rect 363766 150618 394250 150854
rect 394486 150618 424970 150854
rect 425206 150618 455690 150854
rect 455926 150618 486410 150854
rect 486646 150618 517130 150854
rect 517366 150618 547850 150854
rect 548086 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 586302 150854
rect 586538 150618 586622 150854
rect 586858 150618 592650 150854
rect -8726 150586 592650 150618
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 10250 147454
rect 10486 147218 40970 147454
rect 41206 147218 71690 147454
rect 71926 147218 102410 147454
rect 102646 147218 133130 147454
rect 133366 147218 163850 147454
rect 164086 147218 194570 147454
rect 194806 147218 225290 147454
rect 225526 147218 256010 147454
rect 256246 147218 286730 147454
rect 286966 147218 317450 147454
rect 317686 147218 348170 147454
rect 348406 147218 378890 147454
rect 379126 147218 409610 147454
rect 409846 147218 440330 147454
rect 440566 147218 471050 147454
rect 471286 147218 501770 147454
rect 502006 147218 532490 147454
rect 532726 147218 563210 147454
rect 563446 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 10250 147134
rect 10486 146898 40970 147134
rect 41206 146898 71690 147134
rect 71926 146898 102410 147134
rect 102646 146898 133130 147134
rect 133366 146898 163850 147134
rect 164086 146898 194570 147134
rect 194806 146898 225290 147134
rect 225526 146898 256010 147134
rect 256246 146898 286730 147134
rect 286966 146898 317450 147134
rect 317686 146898 348170 147134
rect 348406 146898 378890 147134
rect 379126 146898 409610 147134
rect 409846 146898 440330 147134
rect 440566 146898 471050 147134
rect 471286 146898 501770 147134
rect 502006 146898 532490 147134
rect 532726 146898 563210 147134
rect 563446 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 137494 592650 137526
rect -8726 137258 -8694 137494
rect -8458 137258 -8374 137494
rect -8138 137258 592062 137494
rect 592298 137258 592382 137494
rect 592618 137258 592650 137494
rect -8726 137174 592650 137258
rect -8726 136938 -8694 137174
rect -8458 136938 -8374 137174
rect -8138 136938 592062 137174
rect 592298 136938 592382 137174
rect 592618 136938 592650 137174
rect -8726 136906 592650 136938
rect -8726 133774 592650 133806
rect -8726 133538 -7734 133774
rect -7498 133538 -7414 133774
rect -7178 133538 591102 133774
rect 591338 133538 591422 133774
rect 591658 133538 592650 133774
rect -8726 133454 592650 133538
rect -8726 133218 -7734 133454
rect -7498 133218 -7414 133454
rect -7178 133218 591102 133454
rect 591338 133218 591422 133454
rect 591658 133218 592650 133454
rect -8726 133186 592650 133218
rect -8726 130054 592650 130086
rect -8726 129818 -6774 130054
rect -6538 129818 -6454 130054
rect -6218 129818 590142 130054
rect 590378 129818 590462 130054
rect 590698 129818 592650 130054
rect -8726 129734 592650 129818
rect -8726 129498 -6774 129734
rect -6538 129498 -6454 129734
rect -6218 129498 590142 129734
rect 590378 129498 590462 129734
rect 590698 129498 592650 129734
rect -8726 129466 592650 129498
rect -8726 126334 592650 126366
rect -8726 126098 -5814 126334
rect -5578 126098 -5494 126334
rect -5258 126098 589182 126334
rect 589418 126098 589502 126334
rect 589738 126098 592650 126334
rect -8726 126014 592650 126098
rect -8726 125778 -5814 126014
rect -5578 125778 -5494 126014
rect -5258 125778 589182 126014
rect 589418 125778 589502 126014
rect 589738 125778 592650 126014
rect -8726 125746 592650 125778
rect -8726 122614 592650 122646
rect -8726 122378 -4854 122614
rect -4618 122378 -4534 122614
rect -4298 122378 588222 122614
rect 588458 122378 588542 122614
rect 588778 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -4854 122294
rect -4618 122058 -4534 122294
rect -4298 122058 588222 122294
rect 588458 122058 588542 122294
rect 588778 122058 592650 122294
rect -8726 122026 592650 122058
rect -8726 118894 592650 118926
rect -8726 118658 -3894 118894
rect -3658 118658 -3574 118894
rect -3338 118658 587262 118894
rect 587498 118658 587582 118894
rect 587818 118658 592650 118894
rect -8726 118574 592650 118658
rect -8726 118338 -3894 118574
rect -3658 118338 -3574 118574
rect -3338 118338 587262 118574
rect 587498 118338 587582 118574
rect 587818 118338 592650 118574
rect -8726 118306 592650 118338
rect -8726 115174 592650 115206
rect -8726 114938 -2934 115174
rect -2698 114938 -2614 115174
rect -2378 114938 25610 115174
rect 25846 114938 56330 115174
rect 56566 114938 87050 115174
rect 87286 114938 117770 115174
rect 118006 114938 148490 115174
rect 148726 114938 179210 115174
rect 179446 114938 209930 115174
rect 210166 114938 240650 115174
rect 240886 114938 271370 115174
rect 271606 114938 302090 115174
rect 302326 114938 332810 115174
rect 333046 114938 363530 115174
rect 363766 114938 394250 115174
rect 394486 114938 424970 115174
rect 425206 114938 455690 115174
rect 455926 114938 486410 115174
rect 486646 114938 517130 115174
rect 517366 114938 547850 115174
rect 548086 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 586302 115174
rect 586538 114938 586622 115174
rect 586858 114938 592650 115174
rect -8726 114854 592650 114938
rect -8726 114618 -2934 114854
rect -2698 114618 -2614 114854
rect -2378 114618 25610 114854
rect 25846 114618 56330 114854
rect 56566 114618 87050 114854
rect 87286 114618 117770 114854
rect 118006 114618 148490 114854
rect 148726 114618 179210 114854
rect 179446 114618 209930 114854
rect 210166 114618 240650 114854
rect 240886 114618 271370 114854
rect 271606 114618 302090 114854
rect 302326 114618 332810 114854
rect 333046 114618 363530 114854
rect 363766 114618 394250 114854
rect 394486 114618 424970 114854
rect 425206 114618 455690 114854
rect 455926 114618 486410 114854
rect 486646 114618 517130 114854
rect 517366 114618 547850 114854
rect 548086 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 586302 114854
rect 586538 114618 586622 114854
rect 586858 114618 592650 114854
rect -8726 114586 592650 114618
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 10250 111454
rect 10486 111218 40970 111454
rect 41206 111218 71690 111454
rect 71926 111218 102410 111454
rect 102646 111218 133130 111454
rect 133366 111218 163850 111454
rect 164086 111218 194570 111454
rect 194806 111218 225290 111454
rect 225526 111218 256010 111454
rect 256246 111218 286730 111454
rect 286966 111218 317450 111454
rect 317686 111218 348170 111454
rect 348406 111218 378890 111454
rect 379126 111218 409610 111454
rect 409846 111218 440330 111454
rect 440566 111218 471050 111454
rect 471286 111218 501770 111454
rect 502006 111218 532490 111454
rect 532726 111218 563210 111454
rect 563446 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 10250 111134
rect 10486 110898 40970 111134
rect 41206 110898 71690 111134
rect 71926 110898 102410 111134
rect 102646 110898 133130 111134
rect 133366 110898 163850 111134
rect 164086 110898 194570 111134
rect 194806 110898 225290 111134
rect 225526 110898 256010 111134
rect 256246 110898 286730 111134
rect 286966 110898 317450 111134
rect 317686 110898 348170 111134
rect 348406 110898 378890 111134
rect 379126 110898 409610 111134
rect 409846 110898 440330 111134
rect 440566 110898 471050 111134
rect 471286 110898 501770 111134
rect 502006 110898 532490 111134
rect 532726 110898 563210 111134
rect 563446 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 101494 592650 101526
rect -8726 101258 -8694 101494
rect -8458 101258 -8374 101494
rect -8138 101258 592062 101494
rect 592298 101258 592382 101494
rect 592618 101258 592650 101494
rect -8726 101174 592650 101258
rect -8726 100938 -8694 101174
rect -8458 100938 -8374 101174
rect -8138 100938 592062 101174
rect 592298 100938 592382 101174
rect 592618 100938 592650 101174
rect -8726 100906 592650 100938
rect -8726 97774 592650 97806
rect -8726 97538 -7734 97774
rect -7498 97538 -7414 97774
rect -7178 97538 591102 97774
rect 591338 97538 591422 97774
rect 591658 97538 592650 97774
rect -8726 97454 592650 97538
rect -8726 97218 -7734 97454
rect -7498 97218 -7414 97454
rect -7178 97218 591102 97454
rect 591338 97218 591422 97454
rect 591658 97218 592650 97454
rect -8726 97186 592650 97218
rect -8726 94054 592650 94086
rect -8726 93818 -6774 94054
rect -6538 93818 -6454 94054
rect -6218 93818 590142 94054
rect 590378 93818 590462 94054
rect 590698 93818 592650 94054
rect -8726 93734 592650 93818
rect -8726 93498 -6774 93734
rect -6538 93498 -6454 93734
rect -6218 93498 590142 93734
rect 590378 93498 590462 93734
rect 590698 93498 592650 93734
rect -8726 93466 592650 93498
rect -8726 90334 592650 90366
rect -8726 90098 -5814 90334
rect -5578 90098 -5494 90334
rect -5258 90098 589182 90334
rect 589418 90098 589502 90334
rect 589738 90098 592650 90334
rect -8726 90014 592650 90098
rect -8726 89778 -5814 90014
rect -5578 89778 -5494 90014
rect -5258 89778 589182 90014
rect 589418 89778 589502 90014
rect 589738 89778 592650 90014
rect -8726 89746 592650 89778
rect -8726 86614 592650 86646
rect -8726 86378 -4854 86614
rect -4618 86378 -4534 86614
rect -4298 86378 588222 86614
rect 588458 86378 588542 86614
rect 588778 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -4854 86294
rect -4618 86058 -4534 86294
rect -4298 86058 588222 86294
rect 588458 86058 588542 86294
rect 588778 86058 592650 86294
rect -8726 86026 592650 86058
rect -8726 82894 592650 82926
rect -8726 82658 -3894 82894
rect -3658 82658 -3574 82894
rect -3338 82658 587262 82894
rect 587498 82658 587582 82894
rect 587818 82658 592650 82894
rect -8726 82574 592650 82658
rect -8726 82338 -3894 82574
rect -3658 82338 -3574 82574
rect -3338 82338 587262 82574
rect 587498 82338 587582 82574
rect 587818 82338 592650 82574
rect -8726 82306 592650 82338
rect -8726 79174 592650 79206
rect -8726 78938 -2934 79174
rect -2698 78938 -2614 79174
rect -2378 78938 25610 79174
rect 25846 78938 56330 79174
rect 56566 78938 87050 79174
rect 87286 78938 117770 79174
rect 118006 78938 148490 79174
rect 148726 78938 179210 79174
rect 179446 78938 209930 79174
rect 210166 78938 240650 79174
rect 240886 78938 271370 79174
rect 271606 78938 302090 79174
rect 302326 78938 332810 79174
rect 333046 78938 363530 79174
rect 363766 78938 394250 79174
rect 394486 78938 424970 79174
rect 425206 78938 455690 79174
rect 455926 78938 486410 79174
rect 486646 78938 517130 79174
rect 517366 78938 547850 79174
rect 548086 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 586302 79174
rect 586538 78938 586622 79174
rect 586858 78938 592650 79174
rect -8726 78854 592650 78938
rect -8726 78618 -2934 78854
rect -2698 78618 -2614 78854
rect -2378 78618 25610 78854
rect 25846 78618 56330 78854
rect 56566 78618 87050 78854
rect 87286 78618 117770 78854
rect 118006 78618 148490 78854
rect 148726 78618 179210 78854
rect 179446 78618 209930 78854
rect 210166 78618 240650 78854
rect 240886 78618 271370 78854
rect 271606 78618 302090 78854
rect 302326 78618 332810 78854
rect 333046 78618 363530 78854
rect 363766 78618 394250 78854
rect 394486 78618 424970 78854
rect 425206 78618 455690 78854
rect 455926 78618 486410 78854
rect 486646 78618 517130 78854
rect 517366 78618 547850 78854
rect 548086 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 586302 78854
rect 586538 78618 586622 78854
rect 586858 78618 592650 78854
rect -8726 78586 592650 78618
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 10250 75454
rect 10486 75218 40970 75454
rect 41206 75218 71690 75454
rect 71926 75218 102410 75454
rect 102646 75218 133130 75454
rect 133366 75218 163850 75454
rect 164086 75218 194570 75454
rect 194806 75218 225290 75454
rect 225526 75218 256010 75454
rect 256246 75218 286730 75454
rect 286966 75218 317450 75454
rect 317686 75218 348170 75454
rect 348406 75218 378890 75454
rect 379126 75218 409610 75454
rect 409846 75218 440330 75454
rect 440566 75218 471050 75454
rect 471286 75218 501770 75454
rect 502006 75218 532490 75454
rect 532726 75218 563210 75454
rect 563446 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 10250 75134
rect 10486 74898 40970 75134
rect 41206 74898 71690 75134
rect 71926 74898 102410 75134
rect 102646 74898 133130 75134
rect 133366 74898 163850 75134
rect 164086 74898 194570 75134
rect 194806 74898 225290 75134
rect 225526 74898 256010 75134
rect 256246 74898 286730 75134
rect 286966 74898 317450 75134
rect 317686 74898 348170 75134
rect 348406 74898 378890 75134
rect 379126 74898 409610 75134
rect 409846 74898 440330 75134
rect 440566 74898 471050 75134
rect 471286 74898 501770 75134
rect 502006 74898 532490 75134
rect 532726 74898 563210 75134
rect 563446 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 65494 592650 65526
rect -8726 65258 -8694 65494
rect -8458 65258 -8374 65494
rect -8138 65258 592062 65494
rect 592298 65258 592382 65494
rect 592618 65258 592650 65494
rect -8726 65174 592650 65258
rect -8726 64938 -8694 65174
rect -8458 64938 -8374 65174
rect -8138 64938 592062 65174
rect 592298 64938 592382 65174
rect 592618 64938 592650 65174
rect -8726 64906 592650 64938
rect -8726 61774 592650 61806
rect -8726 61538 -7734 61774
rect -7498 61538 -7414 61774
rect -7178 61538 591102 61774
rect 591338 61538 591422 61774
rect 591658 61538 592650 61774
rect -8726 61454 592650 61538
rect -8726 61218 -7734 61454
rect -7498 61218 -7414 61454
rect -7178 61218 591102 61454
rect 591338 61218 591422 61454
rect 591658 61218 592650 61454
rect -8726 61186 592650 61218
rect -8726 58054 592650 58086
rect -8726 57818 -6774 58054
rect -6538 57818 -6454 58054
rect -6218 57818 590142 58054
rect 590378 57818 590462 58054
rect 590698 57818 592650 58054
rect -8726 57734 592650 57818
rect -8726 57498 -6774 57734
rect -6538 57498 -6454 57734
rect -6218 57498 590142 57734
rect 590378 57498 590462 57734
rect 590698 57498 592650 57734
rect -8726 57466 592650 57498
rect -8726 54334 592650 54366
rect -8726 54098 -5814 54334
rect -5578 54098 -5494 54334
rect -5258 54098 589182 54334
rect 589418 54098 589502 54334
rect 589738 54098 592650 54334
rect -8726 54014 592650 54098
rect -8726 53778 -5814 54014
rect -5578 53778 -5494 54014
rect -5258 53778 589182 54014
rect 589418 53778 589502 54014
rect 589738 53778 592650 54014
rect -8726 53746 592650 53778
rect -8726 50614 592650 50646
rect -8726 50378 -4854 50614
rect -4618 50378 -4534 50614
rect -4298 50378 588222 50614
rect 588458 50378 588542 50614
rect 588778 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -4854 50294
rect -4618 50058 -4534 50294
rect -4298 50058 588222 50294
rect 588458 50058 588542 50294
rect 588778 50058 592650 50294
rect -8726 50026 592650 50058
rect -8726 46894 592650 46926
rect -8726 46658 -3894 46894
rect -3658 46658 -3574 46894
rect -3338 46658 587262 46894
rect 587498 46658 587582 46894
rect 587818 46658 592650 46894
rect -8726 46574 592650 46658
rect -8726 46338 -3894 46574
rect -3658 46338 -3574 46574
rect -3338 46338 587262 46574
rect 587498 46338 587582 46574
rect 587818 46338 592650 46574
rect -8726 46306 592650 46338
rect -8726 43174 592650 43206
rect -8726 42938 -2934 43174
rect -2698 42938 -2614 43174
rect -2378 42938 25610 43174
rect 25846 42938 56330 43174
rect 56566 42938 87050 43174
rect 87286 42938 117770 43174
rect 118006 42938 148490 43174
rect 148726 42938 179210 43174
rect 179446 42938 209930 43174
rect 210166 42938 240650 43174
rect 240886 42938 271370 43174
rect 271606 42938 302090 43174
rect 302326 42938 332810 43174
rect 333046 42938 363530 43174
rect 363766 42938 394250 43174
rect 394486 42938 424970 43174
rect 425206 42938 455690 43174
rect 455926 42938 486410 43174
rect 486646 42938 517130 43174
rect 517366 42938 547850 43174
rect 548086 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 586302 43174
rect 586538 42938 586622 43174
rect 586858 42938 592650 43174
rect -8726 42854 592650 42938
rect -8726 42618 -2934 42854
rect -2698 42618 -2614 42854
rect -2378 42618 25610 42854
rect 25846 42618 56330 42854
rect 56566 42618 87050 42854
rect 87286 42618 117770 42854
rect 118006 42618 148490 42854
rect 148726 42618 179210 42854
rect 179446 42618 209930 42854
rect 210166 42618 240650 42854
rect 240886 42618 271370 42854
rect 271606 42618 302090 42854
rect 302326 42618 332810 42854
rect 333046 42618 363530 42854
rect 363766 42618 394250 42854
rect 394486 42618 424970 42854
rect 425206 42618 455690 42854
rect 455926 42618 486410 42854
rect 486646 42618 517130 42854
rect 517366 42618 547850 42854
rect 548086 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 586302 42854
rect 586538 42618 586622 42854
rect 586858 42618 592650 42854
rect -8726 42586 592650 42618
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 10250 39454
rect 10486 39218 40970 39454
rect 41206 39218 71690 39454
rect 71926 39218 102410 39454
rect 102646 39218 133130 39454
rect 133366 39218 163850 39454
rect 164086 39218 194570 39454
rect 194806 39218 225290 39454
rect 225526 39218 256010 39454
rect 256246 39218 286730 39454
rect 286966 39218 317450 39454
rect 317686 39218 348170 39454
rect 348406 39218 378890 39454
rect 379126 39218 409610 39454
rect 409846 39218 440330 39454
rect 440566 39218 471050 39454
rect 471286 39218 501770 39454
rect 502006 39218 532490 39454
rect 532726 39218 563210 39454
rect 563446 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 10250 39134
rect 10486 38898 40970 39134
rect 41206 38898 71690 39134
rect 71926 38898 102410 39134
rect 102646 38898 133130 39134
rect 133366 38898 163850 39134
rect 164086 38898 194570 39134
rect 194806 38898 225290 39134
rect 225526 38898 256010 39134
rect 256246 38898 286730 39134
rect 286966 38898 317450 39134
rect 317686 38898 348170 39134
rect 348406 38898 378890 39134
rect 379126 38898 409610 39134
rect 409846 38898 440330 39134
rect 440566 38898 471050 39134
rect 471286 38898 501770 39134
rect 502006 38898 532490 39134
rect 532726 38898 563210 39134
rect 563446 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 29494 592650 29526
rect -8726 29258 -8694 29494
rect -8458 29258 -8374 29494
rect -8138 29258 592062 29494
rect 592298 29258 592382 29494
rect 592618 29258 592650 29494
rect -8726 29174 592650 29258
rect -8726 28938 -8694 29174
rect -8458 28938 -8374 29174
rect -8138 28938 592062 29174
rect 592298 28938 592382 29174
rect 592618 28938 592650 29174
rect -8726 28906 592650 28938
rect -8726 25774 592650 25806
rect -8726 25538 -7734 25774
rect -7498 25538 -7414 25774
rect -7178 25538 591102 25774
rect 591338 25538 591422 25774
rect 591658 25538 592650 25774
rect -8726 25454 592650 25538
rect -8726 25218 -7734 25454
rect -7498 25218 -7414 25454
rect -7178 25218 591102 25454
rect 591338 25218 591422 25454
rect 591658 25218 592650 25454
rect -8726 25186 592650 25218
rect -8726 22054 592650 22086
rect -8726 21818 -6774 22054
rect -6538 21818 -6454 22054
rect -6218 21818 590142 22054
rect 590378 21818 590462 22054
rect 590698 21818 592650 22054
rect -8726 21734 592650 21818
rect -8726 21498 -6774 21734
rect -6538 21498 -6454 21734
rect -6218 21498 590142 21734
rect 590378 21498 590462 21734
rect 590698 21498 592650 21734
rect -8726 21466 592650 21498
rect -8726 18334 592650 18366
rect -8726 18098 -5814 18334
rect -5578 18098 -5494 18334
rect -5258 18098 589182 18334
rect 589418 18098 589502 18334
rect 589738 18098 592650 18334
rect -8726 18014 592650 18098
rect -8726 17778 -5814 18014
rect -5578 17778 -5494 18014
rect -5258 17778 589182 18014
rect 589418 17778 589502 18014
rect 589738 17778 592650 18014
rect -8726 17746 592650 17778
rect -8726 14614 592650 14646
rect -8726 14378 -4854 14614
rect -4618 14378 -4534 14614
rect -4298 14378 588222 14614
rect 588458 14378 588542 14614
rect 588778 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -4854 14294
rect -4618 14058 -4534 14294
rect -4298 14058 588222 14294
rect 588458 14058 588542 14294
rect 588778 14058 592650 14294
rect -8726 14026 592650 14058
rect -8726 10894 592650 10926
rect -8726 10658 -3894 10894
rect -3658 10658 -3574 10894
rect -3338 10658 587262 10894
rect 587498 10658 587582 10894
rect 587818 10658 592650 10894
rect -8726 10574 592650 10658
rect -8726 10338 -3894 10574
rect -3658 10338 -3574 10574
rect -3338 10338 587262 10574
rect 587498 10338 587582 10574
rect 587818 10338 592650 10574
rect -8726 10306 592650 10338
rect -8726 7174 592650 7206
rect -8726 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 592650 7174
rect -8726 6854 592650 6938
rect -8726 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 592650 6854
rect -8726 6586 592650 6618
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 41546 -1306
rect 41782 -1542 41866 -1306
rect 42102 -1542 77546 -1306
rect 77782 -1542 77866 -1306
rect 78102 -1542 113546 -1306
rect 113782 -1542 113866 -1306
rect 114102 -1542 149546 -1306
rect 149782 -1542 149866 -1306
rect 150102 -1542 185546 -1306
rect 185782 -1542 185866 -1306
rect 186102 -1542 221546 -1306
rect 221782 -1542 221866 -1306
rect 222102 -1542 257546 -1306
rect 257782 -1542 257866 -1306
rect 258102 -1542 293546 -1306
rect 293782 -1542 293866 -1306
rect 294102 -1542 329546 -1306
rect 329782 -1542 329866 -1306
rect 330102 -1542 365546 -1306
rect 365782 -1542 365866 -1306
rect 366102 -1542 401546 -1306
rect 401782 -1542 401866 -1306
rect 402102 -1542 437546 -1306
rect 437782 -1542 437866 -1306
rect 438102 -1542 473546 -1306
rect 473782 -1542 473866 -1306
rect 474102 -1542 509546 -1306
rect 509782 -1542 509866 -1306
rect 510102 -1542 545546 -1306
rect 545782 -1542 545866 -1306
rect 546102 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 41546 -1626
rect 41782 -1862 41866 -1626
rect 42102 -1862 77546 -1626
rect 77782 -1862 77866 -1626
rect 78102 -1862 113546 -1626
rect 113782 -1862 113866 -1626
rect 114102 -1862 149546 -1626
rect 149782 -1862 149866 -1626
rect 150102 -1862 185546 -1626
rect 185782 -1862 185866 -1626
rect 186102 -1862 221546 -1626
rect 221782 -1862 221866 -1626
rect 222102 -1862 257546 -1626
rect 257782 -1862 257866 -1626
rect 258102 -1862 293546 -1626
rect 293782 -1862 293866 -1626
rect 294102 -1862 329546 -1626
rect 329782 -1862 329866 -1626
rect 330102 -1862 365546 -1626
rect 365782 -1862 365866 -1626
rect 366102 -1862 401546 -1626
rect 401782 -1862 401866 -1626
rect 402102 -1862 437546 -1626
rect 437782 -1862 437866 -1626
rect 438102 -1862 473546 -1626
rect 473782 -1862 473866 -1626
rect 474102 -1862 509546 -1626
rect 509782 -1862 509866 -1626
rect 510102 -1862 545546 -1626
rect 545782 -1862 545866 -1626
rect 546102 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use rift2Wrap  i_Rift2Wrap
timestamp 0
transform 1 0 6000 0 1 6000
box 0 0 570805 686669
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 7375 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 7375 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 7375 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 7375 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 7375 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 7375 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 7375 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 7375 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 7375 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 7375 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 7375 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 7375 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 7375 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 7375 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 7375 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 9234 692105 9854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 45234 692105 45854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 81234 692105 81854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 117234 692460 117854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 153234 692105 153854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 189234 692105 189854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 225234 692460 225854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 261234 692105 261854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 297234 692105 297854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 333234 692105 333854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 369234 692105 369854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 405234 692105 405854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 441234 692105 441854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 692105 477854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 692105 513854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 549234 692105 549854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 10306 592650 10926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 46306 592650 46926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 82306 592650 82926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 118306 592650 118926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 154306 592650 154926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 190306 592650 190926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 226306 592650 226926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 262306 592650 262926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 298306 592650 298926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 334306 592650 334926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 370306 592650 370926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 406306 592650 406926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 442306 592650 442926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 478306 592650 478926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 514306 592650 514926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 550306 592650 550926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 586306 592650 586926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 622306 592650 622926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 658306 592650 658926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 694306 592650 694926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 17746 592650 18366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 53746 592650 54366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 89746 592650 90366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 125746 592650 126366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 161746 592650 162366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 197746 592650 198366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 233746 592650 234366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 269746 592650 270366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 305746 592650 306366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 341746 592650 342366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 377746 592650 378366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 413746 592650 414366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 449746 592650 450366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 485746 592650 486366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 521746 592650 522366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 557746 592650 558366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 593746 592650 594366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 629746 592650 630366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 665746 592650 666366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 25186 592650 25806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 61186 592650 61806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 97186 592650 97806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 133186 592650 133806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 169186 592650 169806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 205186 592650 205806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 241186 592650 241806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 277186 592650 277806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 313186 592650 313806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 349186 592650 349806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 385186 592650 385806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 421186 592650 421806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 457186 592650 457806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 493186 592650 493806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 529186 592650 529806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 565186 592650 565806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 601186 592650 601806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 637186 592650 637806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 673186 592650 673806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 21466 592650 22086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 57466 592650 58086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 93466 592650 94086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 129466 592650 130086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 165466 592650 166086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 201466 592650 202086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 237466 592650 238086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 273466 592650 274086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 309466 592650 310086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 345466 592650 346086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 381466 592650 382086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 417466 592650 418086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 453466 592650 454086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 489466 592650 490086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 525466 592650 526086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 561466 592650 562086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 597466 592650 598086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 633466 592650 634086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 669466 592650 670086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 28906 592650 29526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 64906 592650 65526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 100906 592650 101526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 136906 592650 137526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 172906 592650 173526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 208906 592650 209526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 244906 592650 245526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 280906 592650 281526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 316906 592650 317526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 352906 592650 353526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 388906 592650 389526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 424906 592650 425526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 460906 592650 461526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 496906 592650 497526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 532906 592650 533526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 568906 592650 569526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 604906 592650 605526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 640906 592650 641526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 676906 592650 677526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 5514 -7654 6134 7375 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 41514 -7654 42134 7375 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 77514 -7654 78134 7375 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 113514 -7654 114134 7375 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 149514 -7654 150134 7375 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 185514 -7654 186134 7375 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 221514 -7654 222134 7375 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 257514 -7654 258134 7375 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 293514 -7654 294134 7375 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 329514 -7654 330134 7375 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 365514 -7654 366134 7375 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 401514 -7654 402134 7375 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 437514 -7654 438134 7375 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473514 -7654 474134 7375 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 -7654 510134 7375 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 545514 -7654 546134 7375 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 581514 -7654 582134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 6586 592650 7206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 42586 592650 43206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 78586 592650 79206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 114586 592650 115206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 150586 592650 151206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 186586 592650 187206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 222586 592650 223206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 258586 592650 259206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 294586 592650 295206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 330586 592650 331206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 366586 592650 367206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 402586 592650 403206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 438586 592650 439206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 474586 592650 475206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 510586 592650 511206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 546586 592650 547206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 582586 592650 583206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 618586 592650 619206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 654586 592650 655206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 690586 592650 691206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 12954 692105 13574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 48954 692105 49574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 84954 692105 85574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 120954 692105 121574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 156954 692105 157574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 192954 692105 193574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 228954 692105 229574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 264954 692105 265574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 300954 692105 301574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 336954 692105 337574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 372954 692105 373574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 408954 692460 409574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 444954 692105 445574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 692105 481574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 692460 517574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 552954 692105 553574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 14026 592650 14646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 50026 592650 50646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 86026 592650 86646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 122026 592650 122646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 158026 592650 158646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 194026 592650 194646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 230026 592650 230646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 266026 592650 266646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 302026 592650 302646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 338026 592650 338646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 374026 592650 374646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 410026 592650 410646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 446026 592650 446646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 482026 592650 482646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 518026 592650 518646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 554026 592650 554646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 590026 592650 590646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 626026 592650 626646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 662026 592650 662646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 698026 592650 698646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
rlabel via4 563328 687336 563328 687336 0 vccd1
rlabel metal5 291962 694616 291962 694616 0 vccd2
rlabel metal5 291962 666056 291962 666056 0 vdda1
rlabel metal5 291962 673496 291962 673496 0 vdda2
rlabel metal5 291962 669776 291962 669776 0 vssa1
rlabel metal5 291962 677216 291962 677216 0 vssa2
rlabel via4 547968 655056 547968 655056 0 vssd1
rlabel metal5 291962 698336 291962 698336 0 vssd2
rlabel metal3 583556 284988 583556 284988 0 analog_io[0]
rlabel metal1 443900 699686 443900 699686 0 analog_io[10]
rlabel metal1 379684 699686 379684 699686 0 analog_io[11]
rlabel metal2 314863 692580 314863 692580 0 analog_io[12]
rlabel metal2 251521 692580 251521 692580 0 analog_io[13]
rlabel metal1 187496 695470 187496 695470 0 analog_io[14]
rlabel metal2 121670 698880 121670 698880 0 analog_io[15]
rlabel metal1 59110 700502 59110 700502 0 analog_io[16]
rlabel metal3 1878 697340 1878 697340 0 analog_io[17]
rlabel metal3 4792 633828 4792 633828 0 analog_io[18]
rlabel metal3 4792 583236 4792 583236 0 analog_io[19]
rlabel metal2 579600 336396 579600 336396 0 analog_io[1]
rlabel metal3 1648 540804 1648 540804 0 analog_io[20]
rlabel metal3 1648 488716 1648 488716 0 analog_io[21]
rlabel metal3 4792 431460 4792 431460 0 analog_io[22]
rlabel metal3 1694 384404 1694 384404 0 analog_io[23]
rlabel metal3 1694 332316 1694 332316 0 analog_io[24]
rlabel metal3 3235 280092 3235 280092 0 analog_io[25]
rlabel metal3 4608 229092 4608 229092 0 analog_io[26]
rlabel metal3 1648 175916 1648 175916 0 analog_io[27]
rlabel metal3 1694 123692 1694 123692 0 analog_io[28]
rlabel metal2 579600 388076 579600 388076 0 analog_io[2]
rlabel metal3 581218 444788 581218 444788 0 analog_io[3]
rlabel metal2 579554 494700 579554 494700 0 analog_io[4]
rlabel metal3 581218 551140 581218 551140 0 analog_io[5]
rlabel metal3 581218 604180 581218 604180 0 analog_io[6]
rlabel metal3 581908 657356 581908 657356 0 analog_io[7]
rlabel metal1 571182 695266 571182 695266 0 analog_io[8]
rlabel metal2 504942 693386 504942 693386 0 analog_io[9]
rlabel metal3 581218 6596 581218 6596 0 io_in[0]
rlabel metal2 579554 455396 579554 455396 0 io_in[10]
rlabel metal1 579416 510646 579416 510646 0 io_in[11]
rlabel metal3 581218 564332 581218 564332 0 io_in[12]
rlabel metal3 581218 617508 581218 617508 0 io_in[13]
rlabel via2 578542 659413 578542 659413 0 io_in[14]
rlabel metal2 558946 698299 558946 698299 0 io_in[15]
rlabel metal2 489118 693692 489118 693692 0 io_in[16]
rlabel metal1 427616 699686 427616 699686 0 io_in[17]
rlabel metal2 365010 701634 365010 701634 0 io_in[18]
rlabel metal1 299460 699686 299460 699686 0 io_in[19]
rlabel metal2 579554 49232 579554 49232 0 io_in[1]
rlabel metal2 235697 692580 235697 692580 0 io_in[20]
rlabel metal2 172638 693386 172638 693386 0 io_in[21]
rlabel metal1 107272 700910 107272 700910 0 io_in[22]
rlabel metal1 42366 700366 42366 700366 0 io_in[23]
rlabel metal3 4884 671772 4884 671772 0 io_in[24]
rlabel metal3 4792 621180 4792 621180 0 io_in[25]
rlabel metal3 1878 579972 1878 579972 0 io_in[26]
rlabel metal3 1648 527884 1648 527884 0 io_in[27]
rlabel metal3 4792 469404 4792 469404 0 io_in[28]
rlabel metal3 1648 423572 1648 423572 0 io_in[29]
rlabel metal2 579600 90916 579600 90916 0 io_in[2]
rlabel metal3 1694 371348 1694 371348 0 io_in[30]
rlabel metal3 1694 319260 1694 319260 0 io_in[31]
rlabel metal3 1671 267172 1671 267172 0 io_in[32]
rlabel metal3 1694 214948 1694 214948 0 io_in[33]
rlabel metal3 1694 162860 1694 162860 0 io_in[34]
rlabel metal3 4562 115260 4562 115260 0 io_in[35]
rlabel metal3 4792 77316 4792 77316 0 io_in[36]
rlabel metal3 4792 39372 4792 39372 0 io_in[37]
rlabel metal2 579600 129676 579600 129676 0 io_in[3]
rlabel metal2 579600 168436 579600 168436 0 io_in[4]
rlabel metal2 579600 207196 579600 207196 0 io_in[5]
rlabel metal3 579508 245820 579508 245820 0 io_in[6]
rlabel metal2 579600 297636 579600 297636 0 io_in[7]
rlabel metal2 579600 349316 579600 349316 0 io_in[8]
rlabel metal1 579324 404362 579324 404362 0 io_in[9]
rlabel metal3 581218 33116 581218 33116 0 io_oeb[0]
rlabel metal3 581218 484636 581218 484636 0 io_oeb[10]
rlabel metal2 579554 534004 579554 534004 0 io_oeb[11]
rlabel metal3 581218 590988 581218 590988 0 io_oeb[12]
rlabel metal3 581218 644028 581218 644028 0 io_oeb[13]
rlabel metal3 581218 697204 581218 697204 0 io_oeb[14]
rlabel metal1 523986 695470 523986 695470 0 io_oeb[15]
rlabel metal2 462346 698880 462346 698880 0 io_oeb[16]
rlabel metal1 395600 699686 395600 699686 0 io_oeb[17]
rlabel metal1 331476 699686 331476 699686 0 io_oeb[18]
rlabel metal2 267635 692580 267635 692580 0 io_oeb[19]
rlabel metal3 581218 72964 581218 72964 0 io_oeb[1]
rlabel metal1 202906 695470 202906 695470 0 io_oeb[20]
rlabel metal1 139334 699686 139334 699686 0 io_oeb[21]
rlabel metal2 76130 697578 76130 697578 0 io_oeb[22]
rlabel metal1 11040 700298 11040 700298 0 io_oeb[23]
rlabel metal3 1878 658172 1878 658172 0 io_oeb[24]
rlabel metal3 4792 595884 4792 595884 0 io_oeb[25]
rlabel metal3 4792 545292 4792 545292 0 io_oeb[26]
rlabel metal3 1694 501772 1694 501772 0 io_oeb[27]
rlabel metal3 1694 449548 1694 449548 0 io_oeb[28]
rlabel metal3 1556 397460 1556 397460 0 io_oeb[29]
rlabel via2 578358 116739 578358 116739 0 io_oeb[2]
rlabel metal3 1694 345372 1694 345372 0 io_oeb[30]
rlabel metal3 1694 293148 1694 293148 0 io_oeb[31]
rlabel metal3 1671 241060 1671 241060 0 io_oeb[32]
rlabel metal3 4562 191148 4562 191148 0 io_oeb[33]
rlabel metal3 1694 136748 1694 136748 0 io_oeb[34]
rlabel metal3 1694 84660 1694 84660 0 io_oeb[35]
rlabel metal3 1878 45492 1878 45492 0 io_oeb[36]
rlabel metal3 1878 6460 1878 6460 0 io_oeb[37]
rlabel metal2 579600 155516 579600 155516 0 io_oeb[3]
rlabel metal2 579600 194276 579600 194276 0 io_oeb[4]
rlabel metal3 583556 232764 583556 232764 0 io_oeb[5]
rlabel metal3 579692 272000 579692 272000 0 io_oeb[6]
rlabel metal2 579600 323476 579600 323476 0 io_oeb[7]
rlabel metal2 579554 376788 579554 376788 0 io_oeb[8]
rlabel metal2 579554 429216 579554 429216 0 io_oeb[9]
rlabel metal1 579462 20638 579462 20638 0 io_out[0]
rlabel metal1 579048 471002 579048 471002 0 io_out[10]
rlabel metal3 581218 524484 581218 524484 0 io_out[11]
rlabel metal3 581218 577660 581218 577660 0 io_out[12]
rlabel metal2 578358 620789 578358 620789 0 io_out[13]
rlabel metal2 578358 672639 578358 672639 0 io_out[14]
rlabel metal2 542386 698605 542386 698605 0 io_out[15]
rlabel metal1 475410 695402 475410 695402 0 io_out[16]
rlabel metal2 409945 692580 409945 692580 0 io_out[17]
rlabel metal1 347622 699686 347622 699686 0 io_out[18]
rlabel metal2 283169 692580 283169 692580 0 io_out[19]
rlabel metal1 579554 60690 579554 60690 0 io_out[1]
rlabel metal2 218454 703596 218454 703596 0 io_out[20]
rlabel metal1 155020 695470 155020 695470 0 io_out[21]
rlabel metal1 91126 700706 91126 700706 0 io_out[22]
rlabel metal2 24334 701634 24334 701634 0 io_out[23]
rlabel metal3 4792 659124 4792 659124 0 io_out[24]
rlabel metal3 1878 619140 1878 619140 0 io_out[25]
rlabel metal3 1694 566916 1694 566916 0 io_out[26]
rlabel metal3 4792 507348 4792 507348 0 io_out[27]
rlabel metal3 1648 462604 1648 462604 0 io_out[28]
rlabel metal3 1694 410516 1694 410516 0 io_out[29]
rlabel metal3 581678 99484 581678 99484 0 io_out[2]
rlabel metal3 1694 358428 1694 358428 0 io_out[30]
rlabel metal3 1694 306204 1694 306204 0 io_out[31]
rlabel metal3 3235 254116 3235 254116 0 io_out[32]
rlabel metal3 1694 201892 1694 201892 0 io_out[33]
rlabel metal3 4608 153204 4608 153204 0 io_out[34]
rlabel metal3 1694 97580 1694 97580 0 io_out[35]
rlabel metal3 1694 58548 1694 58548 0 io_out[36]
rlabel metal3 1648 19380 1648 19380 0 io_out[37]
rlabel metal3 582138 139332 582138 139332 0 io_out[3]
rlabel metal3 582046 179180 582046 179180 0 io_out[4]
rlabel metal3 582230 219028 582230 219028 0 io_out[5]
rlabel metal3 580152 258876 580152 258876 0 io_out[6]
rlabel metal2 579600 310556 579600 310556 0 io_out[7]
rlabel metal3 582230 365092 582230 365092 0 io_out[8]
rlabel metal2 579554 416092 579554 416092 0 io_out[9]
rlabel metal2 136206 4668 136206 4668 0 la_data_in[0]
rlabel metal2 467406 4906 467406 4906 0 la_data_in[100]
rlabel metal2 484058 1826 484058 1826 0 la_data_in[101]
rlabel metal2 487646 2098 487646 2098 0 la_data_in[102]
rlabel metal2 477342 5076 477342 5076 0 la_data_in[103]
rlabel metal2 480654 4566 480654 4566 0 la_data_in[104]
rlabel metal2 483966 4838 483966 4838 0 la_data_in[105]
rlabel metal2 487278 4668 487278 4668 0 la_data_in[106]
rlabel metal2 505402 1928 505402 1928 0 la_data_in[107]
rlabel metal2 508898 2234 508898 2234 0 la_data_in[108]
rlabel metal2 497214 5008 497214 5008 0 la_data_in[109]
rlabel metal2 161322 2098 161322 2098 0 la_data_in[10]
rlabel metal2 500802 4709 500802 4709 0 la_data_in[110]
rlabel metal2 503838 4566 503838 4566 0 la_data_in[111]
rlabel metal2 507150 4770 507150 4770 0 la_data_in[112]
rlabel metal2 526654 1588 526654 1588 0 la_data_in[113]
rlabel metal2 513774 5008 513774 5008 0 la_data_in[114]
rlabel metal2 517086 4600 517086 4600 0 la_data_in[115]
rlabel metal2 520398 5042 520398 5042 0 la_data_in[116]
rlabel metal2 526746 3400 526746 3400 0 la_data_in[117]
rlabel metal2 527022 4770 527022 4770 0 la_data_in[118]
rlabel metal2 530334 5008 530334 5008 0 la_data_in[119]
rlabel metal2 172638 4566 172638 4566 0 la_data_in[11]
rlabel metal2 533646 4940 533646 4940 0 la_data_in[120]
rlabel metal2 536958 5042 536958 5042 0 la_data_in[121]
rlabel metal1 544042 3230 544042 3230 0 la_data_in[122]
rlabel metal2 543582 4804 543582 4804 0 la_data_in[123]
rlabel metal2 546894 4634 546894 4634 0 la_data_in[124]
rlabel metal2 550206 5008 550206 5008 0 la_data_in[125]
rlabel metal2 553518 4974 553518 4974 0 la_data_in[126]
rlabel metal2 556830 5042 556830 5042 0 la_data_in[127]
rlabel metal2 175950 5042 175950 5042 0 la_data_in[12]
rlabel metal2 171994 1656 171994 1656 0 la_data_in[13]
rlabel metal2 175490 2064 175490 2064 0 la_data_in[14]
rlabel metal2 179078 2132 179078 2132 0 la_data_in[15]
rlabel metal2 182574 1758 182574 1758 0 la_data_in[16]
rlabel metal2 192510 4532 192510 4532 0 la_data_in[17]
rlabel metal2 195822 5008 195822 5008 0 la_data_in[18]
rlabel metal2 193246 1962 193246 1962 0 la_data_in[19]
rlabel metal2 139518 4770 139518 4770 0 la_data_in[1]
rlabel metal2 196834 1690 196834 1690 0 la_data_in[20]
rlabel metal2 200330 1656 200330 1656 0 la_data_in[21]
rlabel metal2 203918 1758 203918 1758 0 la_data_in[22]
rlabel metal2 212382 4532 212382 4532 0 la_data_in[23]
rlabel metal2 211002 1792 211002 1792 0 la_data_in[24]
rlabel metal2 214498 1656 214498 1656 0 la_data_in[25]
rlabel metal2 218086 2064 218086 2064 0 la_data_in[26]
rlabel metal2 221582 1724 221582 1724 0 la_data_in[27]
rlabel metal2 225170 1656 225170 1656 0 la_data_in[28]
rlabel metal2 232254 4872 232254 4872 0 la_data_in[29]
rlabel metal2 132986 2200 132986 2200 0 la_data_in[2]
rlabel metal2 232254 1656 232254 1656 0 la_data_in[30]
rlabel metal2 235842 1622 235842 1622 0 la_data_in[31]
rlabel metal2 239338 1656 239338 1656 0 la_data_in[32]
rlabel metal2 242926 1622 242926 1622 0 la_data_in[33]
rlabel metal2 248814 4600 248814 4600 0 la_data_in[34]
rlabel metal2 250010 1724 250010 1724 0 la_data_in[35]
rlabel metal2 253506 1690 253506 1690 0 la_data_in[36]
rlabel metal2 257094 1724 257094 1724 0 la_data_in[37]
rlabel metal2 260682 1690 260682 1690 0 la_data_in[38]
rlabel metal2 264178 1724 264178 1724 0 la_data_in[39]
rlabel metal2 136482 2234 136482 2234 0 la_data_in[3]
rlabel metal2 267766 1690 267766 1690 0 la_data_in[40]
rlabel metal2 271262 1724 271262 1724 0 la_data_in[41]
rlabel metal2 274949 204 274949 204 0 la_data_in[42]
rlabel metal2 278346 3203 278346 3203 0 la_data_in[43]
rlabel metal2 281934 3196 281934 3196 0 la_data_in[44]
rlabel metal2 285430 3203 285430 3203 0 la_data_in[45]
rlabel metal2 289018 3203 289018 3203 0 la_data_in[46]
rlabel metal2 292606 1690 292606 1690 0 la_data_in[47]
rlabel metal2 296102 1690 296102 1690 0 la_data_in[48]
rlabel metal2 299690 1758 299690 1758 0 la_data_in[49]
rlabel metal2 140070 2064 140070 2064 0 la_data_in[4]
rlabel metal2 303186 1690 303186 1690 0 la_data_in[50]
rlabel metal2 306774 1724 306774 1724 0 la_data_in[51]
rlabel metal2 310270 1690 310270 1690 0 la_data_in[52]
rlabel metal2 313858 1724 313858 1724 0 la_data_in[53]
rlabel metal2 315054 4566 315054 4566 0 la_data_in[54]
rlabel metal2 320942 1588 320942 1588 0 la_data_in[55]
rlabel metal2 324438 1588 324438 1588 0 la_data_in[56]
rlabel metal2 328026 1724 328026 1724 0 la_data_in[57]
rlabel metal2 331614 1724 331614 1724 0 la_data_in[58]
rlabel metal2 335110 1792 335110 1792 0 la_data_in[59]
rlabel metal2 152766 5042 152766 5042 0 la_data_in[5]
rlabel metal2 334926 4804 334926 4804 0 la_data_in[60]
rlabel metal2 342194 1656 342194 1656 0 la_data_in[61]
rlabel metal2 345782 1758 345782 1758 0 la_data_in[62]
rlabel metal2 349278 1894 349278 1894 0 la_data_in[63]
rlabel metal2 352866 1758 352866 1758 0 la_data_in[64]
rlabel metal2 351486 4498 351486 4498 0 la_data_in[65]
rlabel metal2 359950 1690 359950 1690 0 la_data_in[66]
rlabel metal2 363538 1588 363538 1588 0 la_data_in[67]
rlabel metal2 367034 1656 367034 1656 0 la_data_in[68]
rlabel metal2 370622 1690 370622 1690 0 la_data_in[69]
rlabel metal2 156078 4736 156078 4736 0 la_data_in[6]
rlabel metal2 368046 4498 368046 4498 0 la_data_in[70]
rlabel metal2 371358 4940 371358 4940 0 la_data_in[71]
rlabel metal2 381202 1690 381202 1690 0 la_data_in[72]
rlabel metal2 384790 1656 384790 1656 0 la_data_in[73]
rlabel metal2 388286 2064 388286 2064 0 la_data_in[74]
rlabel metal2 391874 1758 391874 1758 0 la_data_in[75]
rlabel metal2 387918 4532 387918 4532 0 la_data_in[76]
rlabel metal2 391230 4838 391230 4838 0 la_data_in[77]
rlabel metal2 402546 1656 402546 1656 0 la_data_in[78]
rlabel metal2 406042 2098 406042 2098 0 la_data_in[79]
rlabel metal2 159390 5008 159390 5008 0 la_data_in[7]
rlabel metal2 409630 2098 409630 2098 0 la_data_in[80]
rlabel metal2 404478 4770 404478 4770 0 la_data_in[81]
rlabel metal2 407790 5008 407790 5008 0 la_data_in[82]
rlabel metal2 411102 4906 411102 4906 0 la_data_in[83]
rlabel metal2 423798 2030 423798 2030 0 la_data_in[84]
rlabel metal2 427294 2132 427294 2132 0 la_data_in[85]
rlabel metal2 430882 2200 430882 2200 0 la_data_in[86]
rlabel metal2 424350 4940 424350 4940 0 la_data_in[87]
rlabel metal2 427662 4974 427662 4974 0 la_data_in[88]
rlabel metal2 430974 5076 430974 5076 0 la_data_in[89]
rlabel metal2 154238 2200 154238 2200 0 la_data_in[8]
rlabel metal2 445050 2098 445050 2098 0 la_data_in[90]
rlabel metal2 448638 1163 448638 1163 0 la_data_in[91]
rlabel metal2 440910 4634 440910 4634 0 la_data_in[92]
rlabel metal2 444222 4804 444222 4804 0 la_data_in[93]
rlabel metal2 447534 4668 447534 4668 0 la_data_in[94]
rlabel metal2 450846 4872 450846 4872 0 la_data_in[95]
rlabel metal2 466302 1792 466302 1792 0 la_data_in[96]
rlabel metal2 469890 2132 469890 2132 0 la_data_in[97]
rlabel metal2 460782 4770 460782 4770 0 la_data_in[98]
rlabel metal2 464094 5076 464094 5076 0 la_data_in[99]
rlabel metal2 157826 2234 157826 2234 0 la_data_in[9]
rlabel metal2 137310 5008 137310 5008 0 la_data_out[0]
rlabel metal2 468510 4838 468510 4838 0 la_data_out[100]
rlabel metal2 485254 2132 485254 2132 0 la_data_out[101]
rlabel metal2 488842 2030 488842 2030 0 la_data_out[102]
rlabel metal2 478446 5008 478446 5008 0 la_data_out[103]
rlabel metal2 481758 5042 481758 5042 0 la_data_out[104]
rlabel metal2 485070 4600 485070 4600 0 la_data_out[105]
rlabel metal2 488382 4974 488382 4974 0 la_data_out[106]
rlabel metal2 506506 2098 506506 2098 0 la_data_out[107]
rlabel metal2 495006 4872 495006 4872 0 la_data_out[108]
rlabel metal2 498318 5042 498318 5042 0 la_data_out[109]
rlabel metal2 162518 1656 162518 1656 0 la_data_out[10]
rlabel metal2 501906 4675 501906 4675 0 la_data_out[110]
rlabel metal2 504942 4906 504942 4906 0 la_data_out[111]
rlabel metal2 508254 4532 508254 4532 0 la_data_out[112]
rlabel metal2 527850 2030 527850 2030 0 la_data_out[113]
rlabel metal2 514878 4940 514878 4940 0 la_data_out[114]
rlabel metal2 518190 4974 518190 4974 0 la_data_out[115]
rlabel metal2 521502 4753 521502 4753 0 la_data_out[116]
rlabel metal1 526654 3264 526654 3264 0 la_data_out[117]
rlabel metal2 528126 4872 528126 4872 0 la_data_out[118]
rlabel metal2 531438 4566 531438 4566 0 la_data_out[119]
rlabel metal2 173742 4532 173742 4532 0 la_data_out[11]
rlabel metal2 534750 4974 534750 4974 0 la_data_out[120]
rlabel metal2 538062 4685 538062 4685 0 la_data_out[121]
rlabel metal2 541374 4532 541374 4532 0 la_data_out[122]
rlabel metal2 544686 4770 544686 4770 0 la_data_out[123]
rlabel metal2 566858 1724 566858 1724 0 la_data_out[124]
rlabel metal2 551310 4940 551310 4940 0 la_data_out[125]
rlabel metal2 554622 4702 554622 4702 0 la_data_out[126]
rlabel metal2 557934 4906 557934 4906 0 la_data_out[127]
rlabel metal2 177054 4804 177054 4804 0 la_data_out[12]
rlabel metal2 173190 1622 173190 1622 0 la_data_out[13]
rlabel metal2 176686 2200 176686 2200 0 la_data_out[14]
rlabel metal2 180274 2166 180274 2166 0 la_data_out[15]
rlabel metal2 183770 1656 183770 1656 0 la_data_out[16]
rlabel metal2 193614 4770 193614 4770 0 la_data_out[17]
rlabel metal2 190854 1622 190854 1622 0 la_data_out[18]
rlabel metal2 194442 1656 194442 1656 0 la_data_out[19]
rlabel metal2 140622 4702 140622 4702 0 la_data_out[1]
rlabel metal2 197938 2064 197938 2064 0 la_data_out[20]
rlabel metal2 201526 1792 201526 1792 0 la_data_out[21]
rlabel metal2 210174 4566 210174 4566 0 la_data_out[22]
rlabel metal2 213486 4906 213486 4906 0 la_data_out[23]
rlabel metal2 212198 1622 212198 1622 0 la_data_out[24]
rlabel metal2 215694 1724 215694 1724 0 la_data_out[25]
rlabel metal2 219282 1928 219282 1928 0 la_data_out[26]
rlabel metal2 222778 1690 222778 1690 0 la_data_out[27]
rlabel metal2 230046 4566 230046 4566 0 la_data_out[28]
rlabel metal2 229862 1758 229862 1758 0 la_data_out[29]
rlabel metal2 134182 2132 134182 2132 0 la_data_out[2]
rlabel metal2 233450 1690 233450 1690 0 la_data_out[30]
rlabel metal2 237038 1690 237038 1690 0 la_data_out[31]
rlabel metal2 240534 1690 240534 1690 0 la_data_out[32]
rlabel metal2 244122 1690 244122 1690 0 la_data_out[33]
rlabel metal2 249918 4566 249918 4566 0 la_data_out[34]
rlabel metal2 251206 1690 251206 1690 0 la_data_out[35]
rlabel metal2 254702 1724 254702 1724 0 la_data_out[36]
rlabel metal2 258290 1690 258290 1690 0 la_data_out[37]
rlabel metal2 261786 1724 261786 1724 0 la_data_out[38]
rlabel metal2 265374 1622 265374 1622 0 la_data_out[39]
rlabel metal2 137678 2098 137678 2098 0 la_data_out[3]
rlabel metal2 268870 1622 268870 1622 0 la_data_out[40]
rlabel metal2 272603 340 272603 340 0 la_data_out[41]
rlabel metal2 276046 3203 276046 3203 0 la_data_out[42]
rlabel metal2 279542 3203 279542 3203 0 la_data_out[43]
rlabel metal2 283130 3203 283130 3203 0 la_data_out[44]
rlabel metal2 286626 3203 286626 3203 0 la_data_out[45]
rlabel metal2 290023 340 290023 340 0 la_data_out[46]
rlabel metal2 293473 340 293473 340 0 la_data_out[47]
rlabel metal2 296286 4532 296286 4532 0 la_data_out[48]
rlabel metal2 300794 1690 300794 1690 0 la_data_out[49]
rlabel metal2 141266 1928 141266 1928 0 la_data_out[4]
rlabel metal2 304382 1724 304382 1724 0 la_data_out[50]
rlabel metal2 307970 1690 307970 1690 0 la_data_out[51]
rlabel metal2 311466 1588 311466 1588 0 la_data_out[52]
rlabel metal2 315054 1588 315054 1588 0 la_data_out[53]
rlabel metal2 318550 1656 318550 1656 0 la_data_out[54]
rlabel metal2 322138 1724 322138 1724 0 la_data_out[55]
rlabel metal2 325634 1758 325634 1758 0 la_data_out[56]
rlabel metal2 329222 1690 329222 1690 0 la_data_out[57]
rlabel metal2 332718 1622 332718 1622 0 la_data_out[58]
rlabel metal2 332718 4566 332718 4566 0 la_data_out[59]
rlabel metal2 153870 4838 153870 4838 0 la_data_out[5]
rlabel metal2 339894 1690 339894 1690 0 la_data_out[60]
rlabel metal2 343390 1622 343390 1622 0 la_data_out[61]
rlabel metal2 346978 1656 346978 1656 0 la_data_out[62]
rlabel metal2 350474 1724 350474 1724 0 la_data_out[63]
rlabel metal2 354062 1962 354062 1962 0 la_data_out[64]
rlabel metal2 352590 4736 352590 4736 0 la_data_out[65]
rlabel metal2 361146 1622 361146 1622 0 la_data_out[66]
rlabel metal2 364642 1724 364642 1724 0 la_data_out[67]
rlabel metal2 368230 1894 368230 1894 0 la_data_out[68]
rlabel metal2 371726 1826 371726 1826 0 la_data_out[69]
rlabel metal2 157182 4940 157182 4940 0 la_data_out[6]
rlabel metal2 369150 4566 369150 4566 0 la_data_out[70]
rlabel metal2 372462 4770 372462 4770 0 la_data_out[71]
rlabel metal2 382398 1622 382398 1622 0 la_data_out[72]
rlabel metal2 385986 1724 385986 1724 0 la_data_out[73]
rlabel metal2 389482 1962 389482 1962 0 la_data_out[74]
rlabel metal2 393070 1656 393070 1656 0 la_data_out[75]
rlabel metal2 389022 4770 389022 4770 0 la_data_out[76]
rlabel metal2 392334 4702 392334 4702 0 la_data_out[77]
rlabel metal2 403650 1894 403650 1894 0 la_data_out[78]
rlabel metal2 407238 2064 407238 2064 0 la_data_out[79]
rlabel metal2 151846 1690 151846 1690 0 la_data_out[7]
rlabel metal2 410826 1962 410826 1962 0 la_data_out[80]
rlabel metal2 405582 4838 405582 4838 0 la_data_out[81]
rlabel metal2 408894 4974 408894 4974 0 la_data_out[82]
rlabel metal2 412206 4804 412206 4804 0 la_data_out[83]
rlabel metal2 424994 2234 424994 2234 0 la_data_out[84]
rlabel metal2 428490 1894 428490 1894 0 la_data_out[85]
rlabel metal2 422142 4804 422142 4804 0 la_data_out[86]
rlabel metal2 425454 4872 425454 4872 0 la_data_out[87]
rlabel metal2 428766 4770 428766 4770 0 la_data_out[88]
rlabel metal2 442658 2200 442658 2200 0 la_data_out[89]
rlabel metal2 155434 1622 155434 1622 0 la_data_out[8]
rlabel metal2 446246 2064 446246 2064 0 la_data_out[90]
rlabel metal2 449834 1860 449834 1860 0 la_data_out[91]
rlabel metal2 442014 4974 442014 4974 0 la_data_out[92]
rlabel metal2 445326 4736 445326 4736 0 la_data_out[93]
rlabel metal2 448638 5042 448638 5042 0 la_data_out[94]
rlabel metal2 464002 2064 464002 2064 0 la_data_out[95]
rlabel metal2 467498 1860 467498 1860 0 la_data_out[96]
rlabel metal2 458574 4940 458574 4940 0 la_data_out[97]
rlabel metal2 461886 5008 461886 5008 0 la_data_out[98]
rlabel metal2 465198 5042 465198 5042 0 la_data_out[99]
rlabel metal2 158930 1894 158930 1894 0 la_data_out[9]
rlabel metal2 138414 4804 138414 4804 0 la_oenb[0]
rlabel metal2 469614 4702 469614 4702 0 la_oenb[100]
rlabel metal2 486450 1894 486450 1894 0 la_oenb[101]
rlabel metal2 481666 3774 481666 3774 0 la_oenb[102]
rlabel metal2 479550 4804 479550 4804 0 la_oenb[103]
rlabel metal2 482862 4906 482862 4906 0 la_oenb[104]
rlabel metal2 486174 4702 486174 4702 0 la_oenb[105]
rlabel metal2 489486 4736 489486 4736 0 la_oenb[106]
rlabel metal2 507702 1792 507702 1792 0 la_oenb[107]
rlabel metal2 496110 4804 496110 4804 0 la_oenb[108]
rlabel metal2 499422 4838 499422 4838 0 la_oenb[109]
rlabel metal2 171534 4770 171534 4770 0 la_oenb[10]
rlabel metal2 502734 4974 502734 4974 0 la_oenb[110]
rlabel metal2 506046 4736 506046 4736 0 la_oenb[111]
rlabel metal2 525458 1792 525458 1792 0 la_oenb[112]
rlabel metal2 512670 4804 512670 4804 0 la_oenb[113]
rlabel metal2 516074 4709 516074 4709 0 la_oenb[114]
rlabel metal2 519294 4838 519294 4838 0 la_oenb[115]
rlabel metal2 522606 4736 522606 4736 0 la_oenb[116]
rlabel metal2 525918 5076 525918 5076 0 la_oenb[117]
rlabel metal2 546710 2064 546710 2064 0 la_oenb[118]
rlabel metal2 532634 4709 532634 4709 0 la_oenb[119]
rlabel metal2 174846 4906 174846 4906 0 la_oenb[11]
rlabel metal2 535854 4838 535854 4838 0 la_oenb[120]
rlabel metal2 539166 4889 539166 4889 0 la_oenb[121]
rlabel metal2 542478 4736 542478 4736 0 la_oenb[122]
rlabel metal2 545790 4872 545790 4872 0 la_oenb[123]
rlabel metal2 549102 5076 549102 5076 0 la_oenb[124]
rlabel metal2 552414 4821 552414 4821 0 la_oenb[125]
rlabel metal2 555726 4753 555726 4753 0 la_oenb[126]
rlabel metal2 559038 4838 559038 4838 0 la_oenb[127]
rlabel metal2 178158 4736 178158 4736 0 la_oenb[12]
rlabel metal2 174294 2234 174294 2234 0 la_oenb[13]
rlabel metal2 177882 2030 177882 2030 0 la_oenb[14]
rlabel metal2 181470 1792 181470 1792 0 la_oenb[15]
rlabel metal2 191406 4566 191406 4566 0 la_oenb[16]
rlabel metal2 194718 4736 194718 4736 0 la_oenb[17]
rlabel metal2 192050 1758 192050 1758 0 la_oenb[18]
rlabel metal2 195638 1724 195638 1724 0 la_oenb[19]
rlabel metal2 141726 4838 141726 4838 0 la_oenb[1]
rlabel metal2 199134 1894 199134 1894 0 la_oenb[20]
rlabel metal2 202722 1622 202722 1622 0 la_oenb[21]
rlabel metal2 211278 4498 211278 4498 0 la_oenb[22]
rlabel metal2 209806 1588 209806 1588 0 la_oenb[23]
rlabel metal2 213394 1758 213394 1758 0 la_oenb[24]
rlabel metal2 216890 1690 216890 1690 0 la_oenb[25]
rlabel metal2 220478 1656 220478 1656 0 la_oenb[26]
rlabel metal2 223974 1758 223974 1758 0 la_oenb[27]
rlabel metal2 231150 4532 231150 4532 0 la_oenb[28]
rlabel metal2 231058 1724 231058 1724 0 la_oenb[29]
rlabel metal2 135286 1894 135286 1894 0 la_oenb[2]
rlabel metal2 234646 1724 234646 1724 0 la_oenb[30]
rlabel metal2 238142 1724 238142 1724 0 la_oenb[31]
rlabel metal2 241730 1724 241730 1724 0 la_oenb[32]
rlabel metal2 245226 1656 245226 1656 0 la_oenb[33]
rlabel metal2 248814 1690 248814 1690 0 la_oenb[34]
rlabel metal2 252402 1724 252402 1724 0 la_oenb[35]
rlabel metal2 255898 1690 255898 1690 0 la_oenb[36]
rlabel metal2 259486 1724 259486 1724 0 la_oenb[37]
rlabel metal2 262982 1690 262982 1690 0 la_oenb[38]
rlabel metal2 266807 340 266807 340 0 la_oenb[39]
rlabel metal2 138874 2030 138874 2030 0 la_oenb[3]
rlabel metal2 270257 340 270257 340 0 la_oenb[40]
rlabel metal2 273654 3203 273654 3203 0 la_oenb[41]
rlabel metal2 277150 1707 277150 1707 0 la_oenb[42]
rlabel metal2 280738 3203 280738 3203 0 la_oenb[43]
rlabel metal2 284326 1707 284326 1707 0 la_oenb[44]
rlabel metal2 287631 340 287631 340 0 la_oenb[45]
rlabel metal2 291410 1707 291410 1707 0 la_oenb[46]
rlabel metal2 294906 1690 294906 1690 0 la_oenb[47]
rlabel metal2 298494 1690 298494 1690 0 la_oenb[48]
rlabel metal2 301990 1724 301990 1724 0 la_oenb[49]
rlabel metal2 142462 1690 142462 1690 0 la_oenb[4]
rlabel metal2 305578 1690 305578 1690 0 la_oenb[50]
rlabel metal2 309074 1724 309074 1724 0 la_oenb[51]
rlabel metal2 312662 1690 312662 1690 0 la_oenb[52]
rlabel metal2 313950 4532 313950 4532 0 la_oenb[53]
rlabel metal2 319746 1690 319746 1690 0 la_oenb[54]
rlabel metal2 323334 1690 323334 1690 0 la_oenb[55]
rlabel metal2 326830 1656 326830 1656 0 la_oenb[56]
rlabel metal2 330418 1656 330418 1656 0 la_oenb[57]
rlabel metal2 333914 1690 333914 1690 0 la_oenb[58]
rlabel metal2 333822 4498 333822 4498 0 la_oenb[59]
rlabel metal2 154974 4804 154974 4804 0 la_oenb[5]
rlabel metal2 340998 1724 340998 1724 0 la_oenb[60]
rlabel metal2 344586 1690 344586 1690 0 la_oenb[61]
rlabel metal2 348082 1996 348082 1996 0 la_oenb[62]
rlabel metal2 351670 1690 351670 1690 0 la_oenb[63]
rlabel metal2 350382 4464 350382 4464 0 la_oenb[64]
rlabel metal2 353694 4940 353694 4940 0 la_oenb[65]
rlabel metal2 362342 1792 362342 1792 0 la_oenb[66]
rlabel metal2 365838 1758 365838 1758 0 la_oenb[67]
rlabel metal2 369426 1996 369426 1996 0 la_oenb[68]
rlabel metal2 372922 1588 372922 1588 0 la_oenb[69]
rlabel metal2 158286 4974 158286 4974 0 la_oenb[6]
rlabel metal2 370254 4600 370254 4600 0 la_oenb[70]
rlabel metal2 373566 4804 373566 4804 0 la_oenb[71]
rlabel metal2 383594 1758 383594 1758 0 la_oenb[72]
rlabel metal2 387182 1996 387182 1996 0 la_oenb[73]
rlabel metal2 390678 1894 390678 1894 0 la_oenb[74]
rlabel metal2 386814 4566 386814 4566 0 la_oenb[75]
rlabel metal2 390126 4804 390126 4804 0 la_oenb[76]
rlabel metal2 401350 1758 401350 1758 0 la_oenb[77]
rlabel metal2 404846 1690 404846 1690 0 la_oenb[78]
rlabel metal2 408434 2200 408434 2200 0 la_oenb[79]
rlabel metal2 153042 1928 153042 1928 0 la_oenb[7]
rlabel metal2 411930 1724 411930 1724 0 la_oenb[80]
rlabel metal2 406686 4736 406686 4736 0 la_oenb[81]
rlabel metal2 409998 4940 409998 4940 0 la_oenb[82]
rlabel metal2 422602 1928 422602 1928 0 la_oenb[83]
rlabel metal2 426190 2166 426190 2166 0 la_oenb[84]
rlabel metal2 429686 1996 429686 1996 0 la_oenb[85]
rlabel metal2 423246 4906 423246 4906 0 la_oenb[86]
rlabel metal2 426558 5008 426558 5008 0 la_oenb[87]
rlabel metal2 429870 4736 429870 4736 0 la_oenb[88]
rlabel metal2 443854 1962 443854 1962 0 la_oenb[89]
rlabel metal2 156630 1962 156630 1962 0 la_oenb[8]
rlabel metal2 447442 2030 447442 2030 0 la_oenb[90]
rlabel metal2 450938 1928 450938 1928 0 la_oenb[91]
rlabel metal2 443118 4838 443118 4838 0 la_oenb[92]
rlabel metal2 446430 4940 446430 4940 0 la_oenb[93]
rlabel metal2 449742 4600 449742 4600 0 la_oenb[94]
rlabel metal2 465198 1962 465198 1962 0 la_oenb[95]
rlabel metal2 468503 340 468503 340 0 la_oenb[96]
rlabel metal2 459678 4736 459678 4736 0 la_oenb[97]
rlabel metal2 462990 4872 462990 4872 0 la_oenb[98]
rlabel metal2 466302 4804 466302 4804 0 la_oenb[99]
rlabel metal2 160126 2132 160126 2132 0 la_oenb[9]
rlabel metal2 560142 4685 560142 4685 0 user_clock2
rlabel metal2 561246 4736 561246 4736 0 user_irq[0]
rlabel metal2 562350 4804 562350 4804 0 user_irq[1]
rlabel metal2 563454 4770 563454 4770 0 user_irq[2]
rlabel metal2 598 2064 598 2064 0 wb_clk_i
rlabel metal2 1702 2234 1702 2234 0 wb_rst_i
rlabel metal2 2898 1826 2898 1826 0 wbs_ack_o
rlabel metal2 25806 4702 25806 4702 0 wbs_adr_i[0]
rlabel metal2 63342 4600 63342 4600 0 wbs_adr_i[10]
rlabel metal2 51382 1860 51382 1860 0 wbs_adr_i[11]
rlabel metal2 54970 1826 54970 1826 0 wbs_adr_i[12]
rlabel metal2 58466 2166 58466 2166 0 wbs_adr_i[13]
rlabel metal2 62054 2200 62054 2200 0 wbs_adr_i[14]
rlabel metal2 79902 4600 79902 4600 0 wbs_adr_i[15]
rlabel metal2 83214 4532 83214 4532 0 wbs_adr_i[16]
rlabel metal2 72634 1792 72634 1792 0 wbs_adr_i[17]
rlabel metal2 76222 1860 76222 1860 0 wbs_adr_i[18]
rlabel metal2 79718 2064 79718 2064 0 wbs_adr_i[19]
rlabel metal2 12374 1792 12374 1792 0 wbs_adr_i[1]
rlabel metal2 83306 2234 83306 2234 0 wbs_adr_i[20]
rlabel metal2 99774 4770 99774 4770 0 wbs_adr_i[21]
rlabel metal2 103086 4634 103086 4634 0 wbs_adr_i[22]
rlabel metal2 93978 2200 93978 2200 0 wbs_adr_i[23]
rlabel metal2 97474 2234 97474 2234 0 wbs_adr_i[24]
rlabel metal2 101062 2166 101062 2166 0 wbs_adr_i[25]
rlabel metal2 116334 4736 116334 4736 0 wbs_adr_i[26]
rlabel metal2 119646 4974 119646 4974 0 wbs_adr_i[27]
rlabel metal2 111642 1962 111642 1962 0 wbs_adr_i[28]
rlabel metal2 115230 1163 115230 1163 0 wbs_adr_i[29]
rlabel metal2 17066 1928 17066 1928 0 wbs_adr_i[2]
rlabel metal2 118818 1860 118818 1860 0 wbs_adr_i[30]
rlabel metal2 122314 2132 122314 2132 0 wbs_adr_i[31]
rlabel metal2 21850 2234 21850 2234 0 wbs_adr_i[3]
rlabel metal2 43470 4668 43470 4668 0 wbs_adr_i[4]
rlabel metal2 30130 1894 30130 1894 0 wbs_adr_i[5]
rlabel metal2 33626 1860 33626 1860 0 wbs_adr_i[6]
rlabel metal2 37214 1792 37214 1792 0 wbs_adr_i[7]
rlabel metal2 40710 2200 40710 2200 0 wbs_adr_i[8]
rlabel metal2 44298 1724 44298 1724 0 wbs_adr_i[9]
rlabel metal2 4094 1894 4094 1894 0 wbs_cyc_i
rlabel metal2 8786 2098 8786 2098 0 wbs_dat_i[0]
rlabel metal2 64446 4736 64446 4736 0 wbs_dat_i[10]
rlabel metal2 52578 1792 52578 1792 0 wbs_dat_i[11]
rlabel metal2 56074 1996 56074 1996 0 wbs_dat_i[12]
rlabel metal2 59662 1656 59662 1656 0 wbs_dat_i[13]
rlabel metal2 63250 2064 63250 2064 0 wbs_dat_i[14]
rlabel metal2 81006 5076 81006 5076 0 wbs_dat_i[15]
rlabel metal2 70334 1894 70334 1894 0 wbs_dat_i[16]
rlabel metal2 73830 1826 73830 1826 0 wbs_dat_i[17]
rlabel metal2 77418 2200 77418 2200 0 wbs_dat_i[18]
rlabel metal2 80914 1962 80914 1962 0 wbs_dat_i[19]
rlabel metal2 13570 2132 13570 2132 0 wbs_dat_i[1]
rlabel metal2 97566 5008 97566 5008 0 wbs_dat_i[20]
rlabel metal2 100878 4736 100878 4736 0 wbs_dat_i[21]
rlabel metal2 91586 2030 91586 2030 0 wbs_dat_i[22]
rlabel metal2 95174 1860 95174 1860 0 wbs_dat_i[23]
rlabel metal2 98670 1962 98670 1962 0 wbs_dat_i[24]
rlabel metal2 102258 1724 102258 1724 0 wbs_dat_i[25]
rlabel metal2 117438 4770 117438 4770 0 wbs_dat_i[26]
rlabel metal2 120750 4668 120750 4668 0 wbs_dat_i[27]
rlabel metal2 112838 2234 112838 2234 0 wbs_dat_i[28]
rlabel metal2 116426 2098 116426 2098 0 wbs_dat_i[29]
rlabel metal2 18262 1690 18262 1690 0 wbs_dat_i[2]
rlabel metal2 119922 2200 119922 2200 0 wbs_dat_i[30]
rlabel metal2 133998 4906 133998 4906 0 wbs_dat_i[31]
rlabel metal2 23046 2064 23046 2064 0 wbs_dat_i[3]
rlabel metal2 44574 4464 44574 4464 0 wbs_dat_i[4]
rlabel metal2 31326 2030 31326 2030 0 wbs_dat_i[5]
rlabel metal2 34822 1996 34822 1996 0 wbs_dat_i[6]
rlabel metal2 38410 2132 38410 2132 0 wbs_dat_i[7]
rlabel metal2 41906 2064 41906 2064 0 wbs_dat_i[8]
rlabel metal2 45494 1928 45494 1928 0 wbs_dat_i[9]
rlabel metal2 9982 2030 9982 2030 0 wbs_dat_o[0]
rlabel metal2 50186 2030 50186 2030 0 wbs_dat_o[10]
rlabel metal2 53774 2098 53774 2098 0 wbs_dat_o[11]
rlabel metal2 57270 2132 57270 2132 0 wbs_dat_o[12]
rlabel metal2 60858 1724 60858 1724 0 wbs_dat_o[13]
rlabel metal2 64354 1962 64354 1962 0 wbs_dat_o[14]
rlabel metal2 81742 4777 81742 4777 0 wbs_dat_o[15]
rlabel metal2 71530 2098 71530 2098 0 wbs_dat_o[16]
rlabel metal2 75026 2030 75026 2030 0 wbs_dat_o[17]
rlabel metal2 78614 2132 78614 2132 0 wbs_dat_o[18]
rlabel metal2 82110 1996 82110 1996 0 wbs_dat_o[19]
rlabel metal2 14766 1996 14766 1996 0 wbs_dat_o[1]
rlabel metal2 98302 4607 98302 4607 0 wbs_dat_o[20]
rlabel metal2 101982 4940 101982 4940 0 wbs_dat_o[21]
rlabel metal2 92782 2132 92782 2132 0 wbs_dat_o[22]
rlabel metal2 96278 2064 96278 2064 0 wbs_dat_o[23]
rlabel metal2 99866 1996 99866 1996 0 wbs_dat_o[24]
rlabel metal2 103362 2098 103362 2098 0 wbs_dat_o[25]
rlabel metal2 118542 4634 118542 4634 0 wbs_dat_o[26]
rlabel metal2 121854 4906 121854 4906 0 wbs_dat_o[27]
rlabel metal2 114034 1996 114034 1996 0 wbs_dat_o[28]
rlabel metal2 117622 2030 117622 2030 0 wbs_dat_o[29]
rlabel metal2 19458 1724 19458 1724 0 wbs_dat_o[2]
rlabel metal2 121118 1894 121118 1894 0 wbs_dat_o[30]
rlabel metal2 135102 5076 135102 5076 0 wbs_dat_o[31]
rlabel metal2 24242 1758 24242 1758 0 wbs_dat_o[3]
rlabel metal2 28934 1843 28934 1843 0 wbs_dat_o[4]
rlabel metal2 32430 1163 32430 1163 0 wbs_dat_o[5]
rlabel metal2 36018 1588 36018 1588 0 wbs_dat_o[6]
rlabel metal2 39606 2166 39606 2166 0 wbs_dat_o[7]
rlabel metal2 43102 2234 43102 2234 0 wbs_dat_o[8]
rlabel metal2 62238 4804 62238 4804 0 wbs_dat_o[9]
rlabel metal2 11178 1962 11178 1962 0 wbs_sel_i[0]
rlabel metal2 15962 2200 15962 2200 0 wbs_sel_i[1]
rlabel metal2 20654 1911 20654 1911 0 wbs_sel_i[2]
rlabel metal2 25346 1656 25346 1656 0 wbs_sel_i[3]
rlabel metal2 5290 1843 5290 1843 0 wbs_stb_i
rlabel metal2 6486 2166 6486 2166 0 wbs_we_i
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
